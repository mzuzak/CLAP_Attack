// Benchmark "../benchmarks/bench/b14_unroll_syn.v" written by ABC on Fri Sep  3 14:35:13 2021

module b14  ( 
    ADDR_REG_0_, ADDR_REG_10_, ADDR_REG_11_, ADDR_REG_12_, ADDR_REG_13_,
    ADDR_REG_14_, ADDR_REG_15_, ADDR_REG_16_, ADDR_REG_17_, ADDR_REG_18_,
    ADDR_REG_19_, ADDR_REG_1_, ADDR_REG_2_, ADDR_REG_3_, ADDR_REG_4_,
    ADDR_REG_5_, ADDR_REG_6_, ADDR_REG_7_, ADDR_REG_8_, ADDR_REG_9_, B_REG,
    DATAI_0_, DATAI_10_, DATAI_11_, DATAI_12_, DATAI_13_, DATAI_14_,
    DATAI_15_, DATAI_16_, DATAI_17_, DATAI_18_, DATAI_19_, DATAI_1_,
    DATAI_20_, DATAI_21_, DATAI_22_, DATAI_23_, DATAI_24_, DATAI_25_,
    DATAI_26_, DATAI_27_, DATAI_28_, DATAI_29_, DATAI_2_, DATAI_30_,
    DATAI_31_, DATAI_3_, DATAI_4_, DATAI_5_, DATAI_6_, DATAI_7_, DATAI_8_,
    DATAI_9_, DATAO_REG_0_, DATAO_REG_10_, DATAO_REG_11_, DATAO_REG_12_,
    DATAO_REG_13_, DATAO_REG_14_, DATAO_REG_15_, DATAO_REG_16_,
    DATAO_REG_17_, DATAO_REG_18_, DATAO_REG_19_, DATAO_REG_1_,
    DATAO_REG_20_, DATAO_REG_21_, DATAO_REG_22_, DATAO_REG_23_,
    DATAO_REG_24_, DATAO_REG_25_, DATAO_REG_26_, DATAO_REG_27_,
    DATAO_REG_28_, DATAO_REG_29_, DATAO_REG_2_, DATAO_REG_30_,
    DATAO_REG_31_, DATAO_REG_3_, DATAO_REG_4_, DATAO_REG_5_, DATAO_REG_6_,
    DATAO_REG_7_, DATAO_REG_8_, DATAO_REG_9_, D_REG_0_, D_REG_10_,
    D_REG_11_, D_REG_12_, D_REG_13_, D_REG_14_, D_REG_15_, D_REG_16_,
    D_REG_17_, D_REG_18_, D_REG_19_, D_REG_1_, D_REG_20_, D_REG_21_,
    D_REG_22_, D_REG_23_, D_REG_24_, D_REG_25_, D_REG_26_, D_REG_27_,
    D_REG_28_, D_REG_29_, D_REG_2_, D_REG_30_, D_REG_31_, D_REG_3_,
    D_REG_4_, D_REG_5_, D_REG_6_, D_REG_7_, D_REG_8_, D_REG_9_, IR_REG_0_,
    IR_REG_10_, IR_REG_11_, IR_REG_12_, IR_REG_13_, IR_REG_14_, IR_REG_15_,
    IR_REG_16_, IR_REG_17_, IR_REG_18_, IR_REG_19_, IR_REG_1_, IR_REG_20_,
    IR_REG_21_, IR_REG_22_, IR_REG_23_, IR_REG_24_, IR_REG_25_, IR_REG_26_,
    IR_REG_27_, IR_REG_28_, IR_REG_29_, IR_REG_2_, IR_REG_30_, IR_REG_31_,
    IR_REG_3_, IR_REG_4_, IR_REG_5_, IR_REG_6_, IR_REG_7_, IR_REG_8_,
    IR_REG_9_, RD_REG, REG0_REG_0_, REG0_REG_10_, REG0_REG_11_,
    REG0_REG_12_, REG0_REG_13_, REG0_REG_14_, REG0_REG_15_, REG0_REG_16_,
    REG0_REG_17_, REG0_REG_18_, REG0_REG_19_, REG0_REG_1_, REG0_REG_20_,
    REG0_REG_21_, REG0_REG_22_, REG0_REG_23_, REG0_REG_24_, REG0_REG_25_,
    REG0_REG_26_, REG0_REG_27_, REG0_REG_28_, REG0_REG_29_, REG0_REG_2_,
    REG0_REG_30_, REG0_REG_31_, REG0_REG_3_, REG0_REG_4_, REG0_REG_5_,
    REG0_REG_6_, REG0_REG_7_, REG0_REG_8_, REG0_REG_9_, REG1_REG_0_,
    REG1_REG_10_, REG1_REG_11_, REG1_REG_12_, REG1_REG_13_, REG1_REG_14_,
    REG1_REG_15_, REG1_REG_16_, REG1_REG_17_, REG1_REG_18_, REG1_REG_19_,
    REG1_REG_1_, REG1_REG_20_, REG1_REG_21_, REG1_REG_22_, REG1_REG_23_,
    REG1_REG_24_, REG1_REG_25_, REG1_REG_26_, REG1_REG_27_, REG1_REG_28_,
    REG1_REG_29_, REG1_REG_2_, REG1_REG_30_, REG1_REG_31_, REG1_REG_3_,
    REG1_REG_4_, REG1_REG_5_, REG1_REG_6_, REG1_REG_7_, REG1_REG_8_,
    REG1_REG_9_, REG2_REG_0_, REG2_REG_10_, REG2_REG_11_, REG2_REG_12_,
    REG2_REG_13_, REG2_REG_14_, REG2_REG_15_, REG2_REG_16_, REG2_REG_17_,
    REG2_REG_18_, REG2_REG_19_, REG2_REG_1_, REG2_REG_20_, REG2_REG_21_,
    REG2_REG_22_, REG2_REG_23_, REG2_REG_24_, REG2_REG_25_, REG2_REG_26_,
    REG2_REG_27_, REG2_REG_28_, REG2_REG_29_, REG2_REG_2_, REG2_REG_30_,
    REG2_REG_31_, REG2_REG_3_, REG2_REG_4_, REG2_REG_5_, REG2_REG_6_,
    REG2_REG_7_, REG2_REG_8_, REG2_REG_9_, REG3_REG_0_, REG3_REG_10_,
    REG3_REG_11_, REG3_REG_12_, REG3_REG_13_, REG3_REG_14_, REG3_REG_15_,
    REG3_REG_16_, REG3_REG_17_, REG3_REG_18_, REG3_REG_19_, REG3_REG_1_,
    REG3_REG_20_, REG3_REG_21_, REG3_REG_22_, REG3_REG_23_, REG3_REG_24_,
    REG3_REG_25_, REG3_REG_26_, REG3_REG_27_, REG3_REG_28_, REG3_REG_2_,
    REG3_REG_3_, REG3_REG_4_, REG3_REG_5_, REG3_REG_6_, REG3_REG_7_,
    REG3_REG_8_, REG3_REG_9_, STATE_REG, WR_REG,
    n1002, n1006, n1010, n1014, n1018, n1022, n1026, n1030, n1034, n1038,
    n1042, n1046, n1050, n1054, n1058, n1062, n1066, n1070, n1074, n1078,
    n1082, n1086, n1090, n1094, n1098, n1102, n1106, n1110, n1114, n1118,
    n1122, n1126, n1130, n1134, n1138, n1142, n1146, n1150, n1154, n1158,
    n1162, n1166, n1170, n1174, n1178, n1182, n1187, n1192, n1197, n1202,
    n1207, n1212, n1217, n1222, n1227, n1232, n1237, n1242, n1247, n1252,
    n1257, n1262, n1267, n1272, n1277, n1282, n1287, n1292, n1297, n1302,
    n1307, n1312, n1317, n1322, n1327, n1332, n1337, n1341, n174, n179,
    n184, n189, n194, n199, n204, n209, n214, n219, n224, n229, n234, n239,
    n244, n249, n254, n259, n264, n269, n274, n279, n284, n289, n294, n299,
    n304, n309, n314, n319, n324, n329, n334, n339, n344, n349, n354, n359,
    n364, n369, n374, n379, n384, n389, n394, n399, n404, n409, n414, n419,
    n424, n429, n434, n439, n444, n449, n454, n459, n464, n469, n474, n479,
    n484, n489, n494, n499, n504, n509, n514, n519, n524, n529, n534, n539,
    n544, n549, n554, n559, n564, n569, n574, n579, n584, n589, n594, n599,
    n604, n609, n614, n619, n624, n629, n634, n639, n644, n649, n654, n659,
    n664, n669, n674, n679, n684, n689, n694, n699, n704, n709, n714, n719,
    n724, n729, n734, n739, n744, n749, n754, n759, n764, n769, n774, n779,
    n784, n789, n794, n799, n804, n809, n814, n819, n824, n829, n834, n839,
    n844, n849, n854, n859, n864, n869, n874, n879, n884, n889, n894, n899,
    n904, n909, n914, n919, n924, n929, n934, n939, n944, n949, n954, n959,
    n964, n969, n974, n978, n982, n986, n990, n994, n998, keyinput  );
  input  ADDR_REG_0_, ADDR_REG_10_, ADDR_REG_11_, ADDR_REG_12_,
    ADDR_REG_13_, ADDR_REG_14_, ADDR_REG_15_, ADDR_REG_16_, ADDR_REG_17_,
    ADDR_REG_18_, ADDR_REG_19_, ADDR_REG_1_, ADDR_REG_2_, ADDR_REG_3_,
    ADDR_REG_4_, ADDR_REG_5_, ADDR_REG_6_, ADDR_REG_7_, ADDR_REG_8_,
    ADDR_REG_9_, B_REG, DATAI_0_, DATAI_10_, DATAI_11_, DATAI_12_,
    DATAI_13_, DATAI_14_, DATAI_15_, DATAI_16_, DATAI_17_, DATAI_18_,
    DATAI_19_, DATAI_1_, DATAI_20_, DATAI_21_, DATAI_22_, DATAI_23_,
    DATAI_24_, DATAI_25_, DATAI_26_, DATAI_27_, DATAI_28_, DATAI_29_,
    DATAI_2_, DATAI_30_, DATAI_31_, DATAI_3_, DATAI_4_, DATAI_5_, DATAI_6_,
    DATAI_7_, DATAI_8_, DATAI_9_, DATAO_REG_0_, DATAO_REG_10_,
    DATAO_REG_11_, DATAO_REG_12_, DATAO_REG_13_, DATAO_REG_14_,
    DATAO_REG_15_, DATAO_REG_16_, DATAO_REG_17_, DATAO_REG_18_,
    DATAO_REG_19_, DATAO_REG_1_, DATAO_REG_20_, DATAO_REG_21_,
    DATAO_REG_22_, DATAO_REG_23_, DATAO_REG_24_, DATAO_REG_25_,
    DATAO_REG_26_, DATAO_REG_27_, DATAO_REG_28_, DATAO_REG_29_,
    DATAO_REG_2_, DATAO_REG_30_, DATAO_REG_31_, DATAO_REG_3_, DATAO_REG_4_,
    DATAO_REG_5_, DATAO_REG_6_, DATAO_REG_7_, DATAO_REG_8_, DATAO_REG_9_,
    D_REG_0_, D_REG_10_, D_REG_11_, D_REG_12_, D_REG_13_, D_REG_14_,
    D_REG_15_, D_REG_16_, D_REG_17_, D_REG_18_, D_REG_19_, D_REG_1_,
    D_REG_20_, D_REG_21_, D_REG_22_, D_REG_23_, D_REG_24_, D_REG_25_,
    D_REG_26_, D_REG_27_, D_REG_28_, D_REG_29_, D_REG_2_, D_REG_30_,
    D_REG_31_, D_REG_3_, D_REG_4_, D_REG_5_, D_REG_6_, D_REG_7_, D_REG_8_,
    D_REG_9_, IR_REG_0_, IR_REG_10_, IR_REG_11_, IR_REG_12_, IR_REG_13_,
    IR_REG_14_, IR_REG_15_, IR_REG_16_, IR_REG_17_, IR_REG_18_, IR_REG_19_,
    IR_REG_1_, IR_REG_20_, IR_REG_21_, IR_REG_22_, IR_REG_23_, IR_REG_24_,
    IR_REG_25_, IR_REG_26_, IR_REG_27_, IR_REG_28_, IR_REG_29_, IR_REG_2_,
    IR_REG_30_, IR_REG_31_, IR_REG_3_, IR_REG_4_, IR_REG_5_, IR_REG_6_,
    IR_REG_7_, IR_REG_8_, IR_REG_9_, RD_REG, REG0_REG_0_, REG0_REG_10_,
    REG0_REG_11_, REG0_REG_12_, REG0_REG_13_, REG0_REG_14_, REG0_REG_15_,
    REG0_REG_16_, REG0_REG_17_, REG0_REG_18_, REG0_REG_19_, REG0_REG_1_,
    REG0_REG_20_, REG0_REG_21_, REG0_REG_22_, REG0_REG_23_, REG0_REG_24_,
    REG0_REG_25_, REG0_REG_26_, REG0_REG_27_, REG0_REG_28_, REG0_REG_29_,
    REG0_REG_2_, REG0_REG_30_, REG0_REG_31_, REG0_REG_3_, REG0_REG_4_,
    REG0_REG_5_, REG0_REG_6_, REG0_REG_7_, REG0_REG_8_, REG0_REG_9_,
    REG1_REG_0_, REG1_REG_10_, REG1_REG_11_, REG1_REG_12_, REG1_REG_13_,
    REG1_REG_14_, REG1_REG_15_, REG1_REG_16_, REG1_REG_17_, REG1_REG_18_,
    REG1_REG_19_, REG1_REG_1_, REG1_REG_20_, REG1_REG_21_, REG1_REG_22_,
    REG1_REG_23_, REG1_REG_24_, REG1_REG_25_, REG1_REG_26_, REG1_REG_27_,
    REG1_REG_28_, REG1_REG_29_, REG1_REG_2_, REG1_REG_30_, REG1_REG_31_,
    REG1_REG_3_, REG1_REG_4_, REG1_REG_5_, REG1_REG_6_, REG1_REG_7_,
    REG1_REG_8_, REG1_REG_9_, REG2_REG_0_, REG2_REG_10_, REG2_REG_11_,
    REG2_REG_12_, REG2_REG_13_, REG2_REG_14_, REG2_REG_15_, REG2_REG_16_,
    REG2_REG_17_, REG2_REG_18_, REG2_REG_19_, REG2_REG_1_, REG2_REG_20_,
    REG2_REG_21_, REG2_REG_22_, REG2_REG_23_, REG2_REG_24_, REG2_REG_25_,
    REG2_REG_26_, REG2_REG_27_, REG2_REG_28_, REG2_REG_29_, REG2_REG_2_,
    REG2_REG_30_, REG2_REG_31_, REG2_REG_3_, REG2_REG_4_, REG2_REG_5_,
    REG2_REG_6_, REG2_REG_7_, REG2_REG_8_, REG2_REG_9_, REG3_REG_0_,
    REG3_REG_10_, REG3_REG_11_, REG3_REG_12_, REG3_REG_13_, REG3_REG_14_,
    REG3_REG_15_, REG3_REG_16_, REG3_REG_17_, REG3_REG_18_, REG3_REG_19_,
    REG3_REG_1_, REG3_REG_20_, REG3_REG_21_, REG3_REG_22_, REG3_REG_23_,
    REG3_REG_24_, REG3_REG_25_, REG3_REG_26_, REG3_REG_27_, REG3_REG_28_,
    REG3_REG_2_, REG3_REG_3_, REG3_REG_4_, REG3_REG_5_, REG3_REG_6_,
    REG3_REG_7_, REG3_REG_8_, REG3_REG_9_, STATE_REG, WR_REG;
  output n1002, n1006, n1010, n1014, n1018, n1022, n1026, n1030, n1034, n1038,
    n1042, n1046, n1050, n1054, n1058, n1062, n1066, n1070, n1074, n1078,
    n1082, n1086, n1090, n1094, n1098, n1102, n1106, n1110, n1114, n1118,
    n1122, n1126, n1130, n1134, n1138, n1142, n1146, n1150, n1154, n1158,
    n1162, n1166, n1170, n1174, n1178, n1182, n1187, n1192, n1197, n1202,
    n1207, n1212, n1217, n1222, n1227, n1232, n1237, n1242, n1247, n1252,
    n1257, n1262, n1267, n1272, n1277, n1282, n1287, n1292, n1297, n1302,
    n1307, n1312, n1317, n1322, n1327, n1332, n1337, n1341, n174, n179,
    n184, n189, n194, n199, n204, n209, n214, n219, n224, n229, n234, n239,
    n244, n249, n254, n259, n264, n269, n274, n279, n284, n289, n294, n299,
    n304, n309, n314, n319, n324, n329, n334, n339, n344, n349, n354, n359,
    n364, n369, n374, n379, n384, n389, n394, n399, n404, n409, n414, n419,
    n424, n429, n434, n439, n444, n449, n454, n459, n464, n469, n474, n479,
    n484, n489, n494, n499, n504, n509, n514, n519, n524, n529, n534, n539,
    n544, n549, n554, n559, n564, n569, n574, n579, n584, n589, n594, n599,
    n604, n609, n614, n619, n624, n629, n634, n639, n644, n649, n654, n659,
    n664, n669, n674, n679, n684, n689, n694, n699, n704, n709, n714, n719,
    n724, n729, n734, n739, n744, n749, n754, n759, n764, n769, n774, n779,
    n784, n789, n794, n799, n804, n809, n814, n819, n824, n829, n834, n839,
    n844, n849, n854, n859, n864, n869, n874, n879, n884, n889, n894, n899,
    n904, n909, n914, n919, n924, n929, n934, n939, n944, n949, n954, n959,
    n964, n969, n974, n978, n982, n986, n990, n994, n998;
  wire new_n7022_, new_n7031_, new_n7092_, new_n8358_, new_n8909_,
    new_n8064_, new_n8065_, new_n8919_, new_n8920_, new_n8917_, new_n8361_,
    new_n7093_, new_n8938_, new_n8081_, new_n8082_, new_n8364_, new_n8098_,
    new_n8099_, new_n8979_, new_n8984_, new_n8988_, new_n8548_, new_n8367_,
    new_n9001_, new_n9011_, new_n8118_, new_n9016_, new_n9017_, new_n9014_,
    new_n8370_, new_n7094_, new_n9035_, new_n8134_, new_n8135_, new_n8373_,
    new_n9063_, new_n9068_, new_n8153_, new_n9076_, new_n9071_, new_n7095_,
    new_n8376_, new_n9088_, new_n8169_, new_n8170_, new_n9098_, new_n9096_,
    new_n8379_, new_n9131_, new_n7096_, new_n8188_, new_n9136_, new_n9135_,
    new_n9138_, new_n8382_, new_n9153_, new_n8204_, new_n8205_, new_n9163_,
    new_n9100_, new_n9161_, new_n8385_, new_n9183_, new_n9190_, new_n9192_,
    new_n8223_, new_n9195_, new_n8388_, new_n7097_, new_n9206_, new_n8237_,
    new_n8238_, new_n8391_, new_n9226_, new_n9233_, new_n9234_, new_n9239_,
    new_n10578_, new_n8394_, new_n8433_, new_n9254_, new_n8272_,
    new_n8273_, new_n9243_, new_n8295_, new_n8292_, new_n9276_, new_n7098_,
    new_n7032_, new_n10172_, new_n7099_, new_n7100_, new_n9302_,
    new_n9312_, new_n9305_, new_n9314_, new_n9319_, new_n8799_, new_n9303_,
    new_n9350_, new_n9366_, new_n7101_, new_n9381_, new_n9424_, new_n9165_,
    new_n9439_, new_n9454_, new_n9469_, new_n7102_, new_n9483_, new_n9521_,
    new_n10521_, new_n9538_, new_n9549_, new_n9553_, new_n9558_,
    new_n9565_, new_n9579_, new_n9580_, new_n7103_, new_n9593_, new_n9594_,
    new_n9608_, new_n9610_, new_n9623_, new_n9629_, new_n9637_, new_n7774_,
    new_n9638_, new_n9658_, new_n9659_, new_n9673_, new_n9675_, new_n9674_,
    new_n9688_, new_n9581_, new_n7033_, new_n7104_, new_n9708_, new_n9721_,
    new_n9733_, new_n9736_, new_n9738_, new_n9759_, new_n7105_, new_n9773_,
    new_n9787_, new_n9801_, new_n9810_, new_n9813_, new_n9815_, new_n7106_,
    new_n9834_, new_n9836_, new_n9849_, new_n9850_, new_n9864_, new_n9866_,
    new_n7107_, new_n9886_, new_n9897_, new_n9900_, new_n9898_, new_n9923_,
    new_n9924_, new_n9296_, new_n9940_, new_n9943_, new_n9946_, new_n9957_,
    new_n9726_, new_n9968_, new_n9969_, new_n7108_, new_n9983_, new_n9997_,
    new_n9694_, new_n9998_, new_n10004_, new_n10007_, new_n10014_,
    new_n9835_, new_n10022_, new_n8942_, new_n9609_, new_n10030_,
    new_n9926_, new_n10032_, new_n10035_, new_n9740_, new_n10041_,
    new_n10044_, new_n9661_, new_n10053_, new_n7109_, new_n10056_,
    new_n9817_, new_n10062_, new_n10065_, new_n10071_, new_n10049_,
    new_n9970_, new_n9660_, new_n10084_, new_n9925_, new_n7110_,
    new_n10094_, new_n10097_, new_n9547_, new_n9548_, new_n10114_,
    new_n10116_, new_n10127_, new_n10137_, new_n10126_, new_n9842_,
    new_n10069_, new_n10139_, new_n10149_, new_n10156_, new_n10155_,
    new_n10163_, new_n9867_, new_n10171_, new_n10178_, new_n9852_,
    new_n7034_, new_n7111_, new_n10184_, new_n10187_, new_n9640_,
    new_n10194_, new_n10199_, new_n10202_, new_n10207_, new_n10210_,
    new_n9851_, new_n10177_, new_n7112_, new_n10218_, new_n9803_,
    new_n10173_, new_n10227_, new_n10230_, new_n10235_, new_n10240_,
    new_n10243_, new_n10166_, new_n9865_, new_n7113_, new_n10253_,
    new_n9909_, new_n9945_, new_n10152_, new_n10263_, new_n10268_,
    new_n10145_, new_n9595_, new_n10277_, new_n10281_, new_n7114_,
    new_n10291_, new_n10290_, new_n10292_, new_n10297_, new_n10296_,
    new_n10299_, new_n10298_, new_n10306_, new_n10305_, new_n10308_,
    new_n10109_, new_n10307_, new_n10313_, new_n10312_, new_n10314_,
    new_n10315_, new_n10317_, new_n8432_, new_n10322_, new_n8450_,
    new_n7115_, new_n10332_, new_n10370_, new_n10374_, new_n10381_,
    new_n10382_, new_n10388_, new_n10397_, new_n10401_, new_n10369_,
    new_n10367_, new_n8890_, new_n10365_, new_n10363_, new_n10359_,
    new_n10357_, new_n10355_, new_n10350_, new_n10348_, new_n10346_,
    new_n10344_, new_n10340_, new_n7116_, new_n10422_, new_n8650_,
    new_n8564_, new_n8584_, new_n8742_, new_n8762_, new_n8710_,
    new_n10441_, new_n8532_, new_n8467_, new_n8980_, new_n9089_,
    new_n10454_, new_n9228_, new_n9240_, new_n9208_, new_n8880_,
    new_n8911_, new_n8853_, new_n10461_, new_n10463_, new_n7117_,
    new_n8940_, new_n10468_, new_n10470_, new_n8621_, new_n10496_,
    new_n10489_, new_n8586_, new_n8627_, new_n10498_, new_n10504_,
    new_n7035_, new_n10130_, new_n10501_, new_n8910_, new_n10389_,
    new_n10511_, new_n9090_, new_n10516_, new_n10515_, new_n10390_,
    new_n9184_, new_n9207_, new_n7118_, new_n9227_, new_n10522_,
    new_n10510_, new_n10383_, new_n10527_, new_n10539_, new_n10553_,
    new_n10405_, new_n10544_, new_n10556_, new_n7119_, new_n10538_,
    new_n10563_, new_n10566_, new_n10584_, new_n10589_, new_n10592_,
    new_n10590_, new_n10595_, new_n10598_, new_n10601_, new_n7120_,
    new_n10608_, new_n10610_, new_n10613_, new_n10616_, new_n10619_,
    new_n10604_, new_n10625_, new_n10420_, new_n10421_, new_n10334_,
    new_n7731_, new_n10342_, new_n10633_, new_n10352_, new_n10495_,
    new_n10643_, new_n10648_, new_n10651_, new_n10657_, new_n10659_,
    new_n10662_, new_n7121_, new_n10667_, new_n10670_, new_n10668_,
    new_n10672_, new_n10674_, new_n10677_, new_n10679_, new_n10680_,
    new_n9410_, new_n10361_, new_n7122_, new_n10684_, new_n10691_,
    new_n10693_, new_n10697_, new_n10698_, new_n10700_, new_n10702_,
    new_n8895_, new_n7815_, new_n7797_, new_n10730_, new_n7816_,
    new_n7833_, new_n7850_, new_n10758_, new_n7123_, new_n10759_,
    new_n7867_, new_n7884_, new_n10779_, new_n10781_, new_n7901_,
    new_n8985_, new_n10799_, new_n10800_, new_n7935_, new_n7952_,
    new_n10820_, new_n10821_, new_n7969_, new_n7036_, new_n7124_,
    new_n7986_, new_n10840_, new_n10841_, new_n8003_, new_n8020_,
    new_n10861_, new_n10863_, new_n8982_, new_n8037_, new_n10884_,
    new_n8071_, new_n8088_, new_n10902_, new_n10903_, new_n7125_,
    new_n8105_, new_n8124_, new_n10923_, new_n10924_, new_n8141_,
    new_n8159_, new_n7126_, new_n10944_, new_n10946_, new_n8176_,
    new_n10945_, new_n10956_, new_n8194_, new_n8211_, new_n7594_,
    new_n8222_, new_n10983_, new_n8262_, new_n8244_, new_n7127_,
    new_n11015_, new_n11014_, new_n11019_, new_n11021_, new_n11018_,
    new_n11029_, new_n11032_, new_n11034_, new_n11037_, new_n7697_,
    new_n11038_, new_n11049_, new_n11051_, new_n11056_, new_n11054_,
    new_n11058_, new_n11068_, new_n11072_, new_n7128_, new_n11077_,
    new_n11080_, new_n11089_, new_n11087_, new_n11092_, new_n11098_,
    new_n11099_, new_n11105_, new_n11104_, new_n7632_, new_n11107_,
    new_n9873_, new_n11109_, new_n10201_, new_n9272_, new_n9292_,
    new_n11130_, new_n10709_, new_n11137_, new_n10729_, new_n7129_,
    new_n11138_, new_n9681_, new_n11151_, new_n11152_, new_n9396_,
    new_n11153_, new_n11161_, new_n11165_, new_n11170_, new_n7037_,
    new_n7653_, new_n11173_, new_n11183_, new_n11181_, new_n11186_,
    new_n11192_, new_n11193_, new_n11203_, new_n11205_, new_n7130_,
    new_n11210_, new_n11208_, new_n11212_, new_n11220_, new_n11224_,
    new_n11229_, new_n11232_, new_n11241_, new_n7572_, new_n11243_,
    new_n11247_, new_n11245_, new_n11250_, new_n11258_, new_n11262_,
    new_n11267_, new_n11270_, new_n7131_, new_n11279_, new_n11281_,
    new_n11287_, new_n11285_, new_n11289_, new_n11300_, new_n11298_,
    new_n11302_, new_n7766_, new_n7675_, new_n11307_, new_n11310_,
    new_n11290_, new_n11313_, new_n11264_, new_n11316_, new_n11251_,
    new_n11319_, new_n11226_, new_n11322_, new_n7132_, new_n11213_,
    new_n11325_, new_n11188_, new_n11328_, new_n11167_, new_n11331_,
    new_n11094_, new_n11334_, new_n11074_, new_n11337_, new_n7613_,
    new_n11050_, new_n11035_, new_n11344_, new_n11345_, new_n11346_,
    new_n11283_, new_n11347_, new_n11351_, new_n11356_, new_n11362_,
    new_n7133_, new_n11364_, new_n11366_, new_n11370_, new_n11231_,
    new_n11206_, new_n11194_, new_n11382_, new_n11392_, new_n9499_,
    new_n11398_, new_n9724_, new_n11400_, new_n11406_, new_n9516_,
    new_n11079_, new_n11052_, new_n11039_, new_n11420_, new_n11409_,
    new_n11373_, new_n9537_, new_n7134_, new_n11439_, new_n9338_,
    new_n9329_, new_n11457_, new_n11464_, new_n11459_, new_n9536_,
    new_n11471_, new_n9351_, new_n7038_, new_n7135_, new_n9361_,
    new_n9376_, new_n9391_, new_n9405_, new_n9419_, new_n9434_, new_n9449_,
    new_n9464_, new_n9478_, new_n11431_, new_n9794_, new_n9494_,
    new_n9508_, new_n11427_, new_n9530_, new_n9532_, new_n10406_,
    new_n10399_, new_n10391_, new_n10385_, new_n10371_, new_n7136_,
    new_n10372_, new_n10558_, new_n10551_, new_n10572_, new_n10638_,
    new_n10630_, new_n10549_, new_n10546_, new_n10569_, new_n10603_,
    new_n9976_, new_n10628_, new_n10583_, new_n10554_, new_n10542_,
    new_n10565_, new_n10564_, new_n10640_, new_n10641_, new_n10602_,
    new_n10626_, new_n7137_, new_n10482_, new_n10540_, new_n10621_,
    new_n10487_, new_n11410_, new_n7725_, new_n8519_, new_n8670_,
    new_n9139_, new_n8628_, new_n9544_, new_n10229_, new_n10196_,
    new_n10186_, new_n10151_, new_n10034_, new_n10209_, new_n10055_,
    new_n10096_, new_n10006_, new_n9680_, new_n7138_, new_n10426_,
    new_n10536_, new_n10479_, new_n10471_, new_n11341_, new_n11415_,
    new_n11381_, new_n11374_, new_n7591_, new_n7728_, new_n9701_,
    new_n7610_, new_n7629_, new_n7628_, new_n8671_, new_n8833_,
    new_n10413_, new_n8840_, new_n10452_, new_n10396_, new_n10393_,
    new_n7139_, new_n10404_, new_n9155_, new_n9242_, new_n10123_,
    new_n8440_, new_n8445_, new_n8443_, new_n8442_, new_n8473_, new_n8535_,
    new_n9857_, new_n10493_, new_n10433_, new_n8619_, new_n8613_,
    new_n8618_, new_n8623_, new_n10417_, new_n8711_, new_n8713_,
    new_n10414_, new_n9287_, new_n7140_, new_n10503_, new_n8777_,
    new_n8801_, new_n8820_, new_n8821_, new_n8857_, new_n10376_,
    new_n10460_, new_n8921_, new_n8924_, new_n9616_, new_n8941_,
    new_n8967_, new_n9005_, new_n9020_, new_n9091_, new_n9078_, new_n9102_,
    new_n9137_, new_n9167_, new_n10402_, new_n7141_, new_n10284_,
    new_n10283_, new_n9560_, new_n10154_, new_n10165_, new_n10242_,
    new_n9725_, new_n9741_, new_n10157_, new_n10064_, new_n9931_,
    new_n10221_, new_n10174_, new_n10118_, new_n9818_, new_n9647_,
    new_n11117_, new_n10132_, new_n10043_, new_n9902_, new_n9907_,
    new_n7142_, new_n9747_, new_n10260_, new_n9912_, new_n9645_,
    new_n9822_, new_n10220_, new_n9695_, new_n9776_, new_n10336_,
    new_n10337_, new_n9752_, new_n10446_, new_n10447_, new_n10427_,
    new_n10472_, new_n10134_, new_n11136_, new_n11073_, new_n11070_,
    new_n11093_, new_n11171_, new_n7143_, new_n11166_, new_n11187_,
    new_n11184_, new_n11204_, new_n11379_, new_n11225_, new_n11242_,
    new_n11268_, new_n11263_, new_n11280_, new_n11355_, new_n11282_,
    new_n7767_, new_n7587_, new_n7581_, new_n7626_, new_n7621_, new_n7643_,
    new_n7662_, new_n7664_, new_n7683_, new_n7144_, new_n7687_, new_n7706_,
    new_n7708_, new_n8456_, new_n8485_, new_n8549_, new_n8598_,
    new_n10780_, new_n8639_, new_n8660_, new_n11371_, new_n8835_,
    new_n10862_, new_n8867_, new_n8923_, new_n9018_, new_n9021_,
    new_n8255_, new_n11145_, new_n9196_, new_n10278_, new_n7039_,
    new_n7145_, new_n9274_, new_n8418_, new_n8478_, new_n8495_, new_n8471_,
    new_n8541_, new_n8585_, new_n8591_, new_n8609_, new_n8620_, new_n7146_,
    new_n8610_, new_n8617_, new_n8657_, new_n8709_, new_n8719_, new_n8714_,
    new_n8761_, new_n8767_, new_n8788_, new_n8817_, new_n11391_,
    new_n8830_, new_n8856_, new_n8885_, new_n8947_, new_n8964_, new_n8116_,
    new_n9006_, new_n10512_, new_n9036_, new_n9055_, new_n7147_,
    new_n8151_, new_n9060_, new_n9118_, new_n8186_, new_n9172_,
    new_n10523_, new_n8254_, new_n9256_, new_n9285_, new_n9255_,
    new_n11407_, new_n11441_, new_n9582_, new_n9583_, new_n9689_,
    new_n9596_, new_n10271_, new_n9597_, new_n10023_, new_n9612_,
    new_n9611_, new_n7148_, new_n9626_, new_n9641_, new_n9642_, new_n9662_,
    new_n10081_, new_n10050_, new_n9677_, new_n9676_, new_n9684_,
    new_n10170_, new_n7149_, new_n9712_, new_n9723_, new_n9742_,
    new_n9762_, new_n9789_, new_n9804_, new_n9819_, new_n9838_, new_n9837_,
    new_n10015_, new_n9343_, new_n9853_, new_n10215_, new_n10248_,
    new_n9868_, new_n10200_, new_n11110_, new_n11116_, new_n11115_,
    new_n11120_, new_n10121_, new_n7150_, new_n10128_, new_n9746_,
    new_n9899_, new_n9927_, new_n10091_, new_n9971_, new_n10076_,
    new_n9972_, new_n9563_, new_n10000_, new_n9156_, new_n10002_,
    new_n9568_, new_n10070_, new_n10068_, new_n10140_, new_n11446_,
    new_n11451_, new_n10333_, new_n10423_, new_n10466_, new_n7023_,
    new_n9120_, new_n7151_, new_n10467_, new_n10734_, new_n10733_,
    new_n10744_, new_n10743_, new_n10765_, new_n10764_, new_n10794_,
    new_n10793_, new_n10826_, new_n8696_, new_n10825_, new_n10855_,
    new_n10854_, new_n10888_, new_n10887_, new_n10896_, new_n10895_,
    new_n10909_, new_n10908_, new_n10917_, new_n7152_, new_n10916_,
    new_n10930_, new_n10929_, new_n10938_, new_n10937_, new_n10951_,
    new_n10950_, new_n10970_, new_n10969_, new_n10712_, new_n9748_,
    new_n10995_, new_n10994_, new_n11003_, new_n11002_, new_n10713_,
    new_n11411_, new_n11163_, new_n11385_, new_n11222_, new_n11375_,
    new_n7153_, new_n11260_, new_n11358_, new_n7603_, new_n10694_,
    new_n7701_, new_n10757_, new_n10778_, new_n7929_, new_n10819_,
    new_n7946_, new_n9648_, new_n10839_, new_n10860_, new_n8863_,
    new_n8054_, new_n10901_, new_n10922_, new_n10943_, new_n8300_,
    new_n8256_, new_n9275_, new_n7154_, new_n8426_, new_n8425_, new_n8451_,
    new_n8496_, new_n8815_, new_n8962_, new_n8998_, new_n9053_, new_n9116_,
    new_n9150_, new_n10455_, new_n9283_, new_n8290_, new_n10318_,
    new_n11460_, new_n11465_, new_n9555_, new_n9737_, new_n9551_,
    new_n9814_, new_n9937_, new_n7155_, new_n9939_, new_n10707_,
    new_n10723_, new_n8454_, new_n8483_, new_n10751_, new_n8552_,
    new_n10772_, new_n10785_, new_n8637_, new_n7156_, new_n10804_,
    new_n10813_, new_n8729_, new_n10833_, new_n10846_, new_n8805_,
    new_n10867_, new_n10875_, new_n8927_, new_n8928_, new_n7040_,
    new_n9711_, new_n8952_, new_n9024_, new_n9025_, new_n9043_, new_n9075_,
    new_n10959_, new_n9173_, new_n10977_, new_n10986_, new_n9216_,
    new_n7157_, new_n10442_, new_n11132_, new_n7580_, new_n11016_,
    new_n11421_, new_n7589_, new_n11401_, new_n11095_, new_n11060_,
    new_n11189_, new_n9911_, new_n11304_, new_n11303_, new_n10663_,
    new_n7645_, new_n10685_, new_n7690_, new_n11434_, new_n7782_,
    new_n7803_, new_n7823_, new_n7158_, new_n7840_, new_n7857_, new_n7874_,
    new_n7891_, new_n7908_, new_n7925_, new_n7942_, new_n7959_, new_n7976_,
    new_n7993_, new_n7159_, new_n8015_, new_n8010_, new_n8032_, new_n8027_,
    new_n8044_, new_n8066_, new_n8061_, new_n8078_, new_n8095_, new_n8112_,
    new_n8726_, new_n8136_, new_n8131_, new_n8148_, new_n8166_, new_n8189_,
    new_n8183_, new_n8201_, new_n7793_, new_n8234_, new_n8251_, new_n7160_,
    new_n8269_, new_n8297_, new_n7790_, new_n8422_, new_n8462_, new_n8459_,
    new_n8474_, new_n8488_, new_n8504_, new_n8527_, new_n7161_, new_n8524_,
    new_n8537_, new_n8559_, new_n8556_, new_n8565_, new_n8578_, new_n8575_,
    new_n8587_, new_n8604_, new_n8601_, new_n9320_, new_n8630_, new_n8645_,
    new_n8642_, new_n8653_, new_n8680_, new_n8677_, new_n8686_, new_n8704_,
    new_n8701_, new_n8715_, new_n7162_, new_n8737_, new_n8734_, new_n8743_,
    new_n8756_, new_n8753_, new_n8763_, new_n8783_, new_n8780_, new_n8790_,
    new_n8811_, new_n9057_, new_n9470_, new_n8808_, new_n8826_, new_n8848_,
    new_n8845_, new_n8858_, new_n8875_, new_n8872_, new_n8881_, new_n8905_,
    new_n8902_, new_n7163_, new_n8912_, new_n8934_, new_n8931_, new_n8943_,
    new_n8958_, new_n8955_, new_n8973_, new_n8995_, new_n8992_, new_n9007_,
    new_n9382_, new_n9031_, new_n9028_, new_n9037_, new_n9049_, new_n9046_,
    new_n9064_, new_n9084_, new_n9081_, new_n9092_, new_n9112_, new_n7164_,
    new_n9109_, new_n9127_, new_n9147_, new_n9144_, new_n9157_, new_n9179_,
    new_n9176_, new_n9186_, new_n9202_, new_n9199_, new_n9367_, new_n9209_,
    new_n9222_, new_n9219_, new_n9229_, new_n9250_, new_n9247_, new_n9257_,
    new_n8398_, new_n9267_, new_n9336_, new_n7165_, new_n9389_, new_n9403_,
    new_n9485_, new_n9506_, new_n9523_, new_n9543_, new_n9541_, new_n9571_,
    new_n9569_, new_n9575_, new_n8669_, new_n9586_, new_n9584_, new_n9589_,
    new_n9600_, new_n9598_, new_n9604_, new_n9615_, new_n9613_, new_n9619_,
    new_n9627_, new_n7166_, new_n9633_, new_n9651_, new_n9649_, new_n9654_,
    new_n9665_, new_n9663_, new_n9669_, new_n9700_, new_n9698_, new_n9704_,
    new_n8697_, new_n9713_, new_n9717_, new_n9729_, new_n9727_, new_n9751_,
    new_n9749_, new_n9755_, new_n9765_, new_n9763_, new_n9769_, new_n7167_,
    new_n9780_, new_n9778_, new_n9783_, new_n9793_, new_n9791_, new_n9797_,
    new_n9807_, new_n9805_, new_n9826_, new_n9824_, new_n7041_, new_n7168_,
    new_n9830_, new_n9841_, new_n9839_, new_n9845_, new_n9856_, new_n9854_,
    new_n9860_, new_n9869_, new_n9878_, new_n9876_, new_n10159_,
    new_n9882_, new_n9890_, new_n9888_, new_n9893_, new_n9915_, new_n9913_,
    new_n9919_, new_n9930_, new_n9928_, new_n9934_, new_n7169_, new_n9949_,
    new_n9953_, new_n9961_, new_n9959_, new_n9964_, new_n9975_, new_n9973_,
    new_n9979_, new_n9989_, new_n9987_, new_n9425_, new_n9993_,
    new_n10104_, new_n10102_, new_n10110_, new_n10329_, new_n8419_,
    new_n8429_, new_n10717_, new_n10724_, new_n10752_, new_n7170_,
    new_n10773_, new_n10786_, new_n10805_, new_n10814_, new_n10834_,
    new_n10847_, new_n10868_, new_n10876_, new_n10960_, new_n10978_,
    new_n9440_, new_n10987_, new_n11133_, new_n11011_, new_n11028_,
    new_n11025_, new_n11042_, new_n11040_, new_n11061_, new_n11083_,
    new_n11081_, new_n7171_, new_n11154_, new_n11174_, new_n11195_,
    new_n11214_, new_n11233_, new_n11252_, new_n11271_, new_n11291_,
    new_n7570_, new_n7592_, new_n9455_, new_n7611_, new_n7630_, new_n7651_,
    new_n7673_, new_n7695_, new_n7768_, new_n7776_, new_n7784_, new_n7791_,
    new_n7810_, new_n7172_, new_n7811_, new_n7829_, new_n7830_, new_n7846_,
    new_n7847_, new_n7863_, new_n7864_, new_n7880_, new_n7881_, new_n7897_,
    new_n7173_, new_n7898_, new_n7914_, new_n7915_, new_n7931_, new_n7932_,
    new_n7948_, new_n7949_, new_n7965_, new_n7966_, new_n7982_, new_n8824_,
    new_n7174_, new_n7983_, new_n7999_, new_n8000_, new_n8016_, new_n8017_,
    new_n8033_, new_n8034_, new_n8050_, new_n8051_, new_n8067_, new_n7175_,
    new_n8068_, new_n8084_, new_n8085_, new_n8101_, new_n8102_, new_n8120_,
    new_n8121_, new_n8137_, new_n8138_, new_n8155_, new_n7176_, new_n8156_,
    new_n8172_, new_n8173_, new_n8190_, new_n8191_, new_n8207_, new_n8208_,
    new_n8224_, new_n8225_, new_n8218_, new_n8518_, new_n8240_, new_n8241_,
    new_n8258_, new_n8259_, new_n8275_, new_n8276_, new_n8282_, new_n8293_,
    new_n8303_, new_n8307_, new_n7177_, new_n8423_, new_n8460_, new_n8489_,
    new_n8525_, new_n8557_, new_n8576_, new_n8602_, new_n8643_, new_n8678_,
    new_n8702_, new_n8513_, new_n8735_, new_n8754_, new_n8781_, new_n8809_,
    new_n8846_, new_n8873_, new_n8903_, new_n8932_, new_n8956_, new_n8993_,
    new_n7178_, new_n9029_, new_n9047_, new_n9082_, new_n9110_, new_n9145_,
    new_n9177_, new_n9200_, new_n9220_, new_n9248_, new_n8397_, new_n8666_,
    new_n9263_, new_n9309_, new_n9325_, new_n9333_, new_n9347_, new_n9356_,
    new_n9371_, new_n9386_, new_n9395_, new_n9400_, new_n7179_, new_n9409_,
    new_n9414_, new_n9429_, new_n9444_, new_n9459_, new_n9474_, new_n9489_,
    new_n9503_, new_n9512_, new_n9527_, new_n8896_, new_n9570_, new_n9599_,
    new_n9628_, new_n9664_, new_n9714_, new_n9728_, new_n9764_, new_n9825_,
    new_n9870_, new_n9877_, new_n7042_, new_n7180_, new_n9914_, new_n9950_,
    new_n9988_, new_n11041_, new_n11062_, new_n11155_, new_n11175_,
    new_n11196_, new_n11215_, new_n11234_, new_n7181_, new_n11253_,
    new_n11272_, new_n11292_, new_n7571_, new_n7593_, new_n7612_,
    new_n7631_, new_n7652_, new_n7674_, new_n7696_, new_n8986_, new_n7769_,
    new_n7777_, new_n7785_, new_n8283_, new_n9306_, new_n9315_, new_n9322_,
    new_n9330_, new_n9339_, new_n9344_, new_n7182_, new_n9353_, new_n9362_,
    new_n9368_, new_n9377_, new_n9383_, new_n9392_, new_n9397_, new_n9406_,
    new_n9411_, new_n9420_, new_n7183_, new_n9426_, new_n9435_, new_n9441_,
    new_n9450_, new_n9456_, new_n9465_, new_n9471_, new_n9479_, new_n9486_,
    new_n9495_, new_n7184_, new_n9500_, new_n9509_, new_n9517_, new_n9524_,
    new_n8750_, new_n8100_, new_n8774_, new_n8521_, new_n8869_, new_n8553_,
    new_n8221_, new_n8674_, new_n8841_, new_n9106_, new_n9171_, new_n8728_,
    new_n8206_, new_n7964_, new_n8596_, new_n8257_, new_n8154_, new_n7185_,
    new_n8119_, new_n10586_, new_n9278_, new_n11036_, new_n11417_,
    new_n9166_, new_n8794_, new_n8916_, new_n8152_, new_n11066_,
    new_n7186_, new_n10531_, new_n10033_, new_n10054_, new_n10095_,
    new_n10185_, new_n10195_, new_n10241_, new_n10164_, new_n10042_,
    new_n10005_, new_n7187_, new_n10063_, new_n10208_, new_n10228_,
    new_n10150_, new_n10219_, new_n11114_, new_n7981_, new_n8239_,
    new_n10703_, new_n7722_, new_n8971_, new_n10158_, new_n9265_,
    new_n8731_, new_n8690_, new_n9300_, new_n8551_, new_n8572_,
    new_n11017_, new_n10596_, new_n7689_, new_n9775_, new_n7188_,
    new_n8444_, new_n8891_, new_n9133_, new_n9944_, new_n10649_,
    new_n10611_, new_n7646_, new_n7609_, new_n8468_, new_n10378_,
    new_n7189_, new_n7819_, new_n7836_, new_n7853_, new_n7870_, new_n7887_,
    new_n7904_, new_n7921_, new_n7938_, new_n7955_, new_n7972_, new_n7190_,
    new_n7989_, new_n8006_, new_n8023_, new_n8040_, new_n8057_, new_n8074_,
    new_n8091_, new_n8108_, new_n8127_, new_n8144_, new_n7191_, new_n8162_,
    new_n8179_, new_n8197_, new_n8214_, new_n8230_, new_n8247_, new_n8265_,
    new_n8281_, new_n8667_, new_n8981_, new_n7192_, new_n7657_, new_n8304_,
    new_n8115_, new_n9554_, new_n8171_, new_n7998_, new_n9235_, new_n8083_,
    new_n8049_, new_n9293_, new_n7193_, new_n8274_, new_n7798_, new_n8291_,
    new_n10122_, new_n11159_, new_n11106_, new_n8536_, new_n9948_,
    new_n9905_, new_n9821_, new_n7194_, new_n9745_, new_n9567_, new_n9986_,
    new_n11090_, new_n11248_, new_n8968_, new_n10652_, new_n8472_,
    new_n10319_, new_n8899_, new_n7195_, new_n9432_, new_n9447_,
    new_n9417_, new_n10119_, new_n10138_, new_n8969_, new_n8629_,
    new_n8854_, new_n10411_, new_n9646_, new_n10279_, new_n10415_,
    new_n9492_, new_n10375_, new_n8615_, new_n8512_, new_n7617_,
    new_n7576_, new_n7605_, new_n10614_, new_n10617_, new_n7043_,
    new_n7196_, new_n10464_, new_n8413_, new_n7772_, new_n8747_,
    new_n8862_, new_n8117_, new_n8187_, new_n11179_, new_n8822_,
    new_n7738_, new_n7197_, new_n10416_, new_n8989_, new_n8502_,
    new_n9126_, new_n8614_, new_n8399_, new_n9282_, new_n10635_,
    new_n9685_, new_n8407_, new_n7198_, new_n9122_, new_n9059_, new_n9359_,
    new_n9374_, new_n9462_, new_n7739_, new_n10593_, new_n7574_,
    new_n4556_, new_n7596_, new_n9632_, new_n4557_, new_n7615_, new_n4558_,
    new_n7634_, new_n4559_, new_n7655_, new_n4560_, new_n7677_, new_n4561_,
    new_n7699_, new_n7199_, new_n4562_, new_n7713_, new_n4563_, new_n7716_,
    new_n4564_, new_n7719_, new_n4565_, new_n7724_, new_n4566_, new_n7730_,
    new_n7200_, new_n4567_, new_n7742_, new_n4568_, new_n7745_, new_n4569_,
    new_n7748_, new_n4570_, new_n7751_, new_n4571_, new_n7755_, new_n7201_,
    new_n4572_, new_n7759_, new_n4573_, new_n7763_, new_n4574_, new_n7770_,
    new_n4575_, new_n7773_, new_n4576_, new_n7778_, new_n7202_, new_n4577_,
    new_n7780_, new_n4578_, new_n7795_, new_n4579_, new_n7804_, new_n4580_,
    new_n7812_, new_n4581_, new_n7817_, new_n7203_, new_n4582_, new_n7824_,
    new_n4583_, new_n7831_, new_n4584_, new_n7834_, new_n4585_, new_n7841_,
    new_n4586_, new_n7848_, new_n7204_, new_n4587_, new_n7851_, new_n4588_,
    new_n7858_, new_n4589_, new_n7865_, new_n4590_, new_n7868_, new_n4591_,
    new_n7875_, new_n7044_, new_n7205_, new_n4592_, new_n7882_, new_n4593_,
    new_n7885_, new_n4594_, new_n7892_, new_n4595_, new_n7899_, new_n4596_,
    new_n7902_, new_n7206_, new_n4597_, new_n7909_, new_n4598_, new_n7916_,
    new_n4599_, new_n7919_, new_n4600_, new_n7926_, new_n4601_, new_n7933_,
    new_n7733_, new_n4602_, new_n7936_, new_n4603_, new_n7943_, new_n4604_,
    new_n7950_, new_n4605_, new_n7953_, new_n4606_, new_n7960_, new_n7207_,
    new_n4607_, new_n7967_, new_n4608_, new_n7970_, new_n4609_, new_n7977_,
    new_n4610_, new_n7984_, new_n4611_, new_n7987_, new_n7208_, new_n4612_,
    new_n7994_, new_n4613_, new_n8001_, new_n4614_, new_n8004_, new_n4615_,
    new_n8011_, new_n4616_, new_n8018_, new_n11357_, new_n4617_,
    new_n8021_, new_n4618_, new_n8028_, new_n4619_, new_n8035_, new_n4620_,
    new_n8038_, new_n4621_, new_n8045_, new_n7209_, new_n4622_, new_n8052_,
    new_n4623_, new_n8055_, new_n4624_, new_n8062_, new_n4625_, new_n8069_,
    new_n4626_, new_n8072_, new_n11393_, new_n4627_, new_n8079_,
    new_n4628_, new_n8086_, new_n4629_, new_n8089_, new_n4630_, new_n8096_,
    new_n4631_, new_n8103_, new_n7210_, new_n4632_, new_n8106_, new_n4633_,
    new_n8113_, new_n4634_, new_n8122_, new_n4635_, new_n8125_, new_n4636_,
    new_n8132_, new_n8972_, new_n4637_, new_n8139_, new_n4638_, new_n8142_,
    new_n4639_, new_n8149_, new_n4640_, new_n8157_, new_n4641_, new_n8160_,
    new_n7045_, new_n7211_, new_n4642_, new_n8167_, new_n4643_, new_n8174_,
    new_n4644_, new_n8177_, new_n4645_, new_n8184_, new_n4646_, new_n8192_,
    new_n9121_, new_n4647_, new_n8195_, new_n4648_, new_n8202_, new_n4649_,
    new_n8209_, new_n4650_, new_n8212_, new_n4651_, new_n8219_, new_n7212_,
    new_n4652_, new_n8226_, new_n4653_, new_n8228_, new_n4654_, new_n8235_,
    new_n4655_, new_n8242_, new_n4656_, new_n8245_, new_n10801_,
    new_n4657_, new_n8252_, new_n4658_, new_n8260_, new_n4659_, new_n8263_,
    new_n4660_, new_n8270_, new_n4661_, new_n8277_, new_n7213_, new_n4662_,
    new_n8279_, new_n4663_, new_n8299_, new_n4664_, new_n8296_, new_n4665_,
    new_n8410_, new_n4666_, new_n8430_, new_n10440_, new_n4667_,
    new_n8427_, new_n4668_, new_n8441_, new_n4669_, new_n8446_, new_n4670_,
    new_n8434_, new_n4671_, new_n8447_, new_n7214_, new_n4672_, new_n8452_,
    new_n4673_, new_n8464_, new_n4674_, new_n8476_, new_n4675_, new_n8497_,
    new_n4676_, new_n8499_, new_n7215_, new_n4677_, new_n8506_, new_n4678_,
    new_n8509_, new_n4679_, new_n8520_, new_n4680_, new_n8529_, new_n4681_,
    new_n8539_, new_n7216_, new_n4682_, new_n8561_, new_n4683_, new_n8567_,
    new_n4684_, new_n8580_, new_n4685_, new_n8589_, new_n4686_, new_n8594_,
    new_n7217_, new_n4687_, new_n8606_, new_n4688_, new_n8632_, new_n4689_,
    new_n8647_, new_n4690_, new_n8655_, new_n4691_, new_n8662_, new_n7024_,
    new_n7046_, new_n7218_, new_n4692_, new_n8682_, new_n4693_, new_n8688_,
    new_n4694_, new_n8691_, new_n4695_, new_n8695_, new_n4696_, new_n8706_,
    new_n7219_, new_n4697_, new_n8720_, new_n4698_, new_n8717_, new_n4699_,
    new_n8722_, new_n4700_, new_n8739_, new_n4701_, new_n8745_, new_n7220_,
    new_n4702_, new_n8758_, new_n4703_, new_n8768_, new_n4704_, new_n8765_,
    new_n4705_, new_n8785_, new_n4706_, new_n8792_, new_n7221_, new_n4707_,
    new_n8802_, new_n4708_, new_n8804_, new_n4709_, new_n8816_, new_n4710_,
    new_n8813_, new_n4711_, new_n8831_, new_n7222_, new_n4712_, new_n8828_,
    new_n4713_, new_n8836_, new_n4714_, new_n8850_, new_n4715_, new_n8860_,
    new_n4716_, new_n8877_, new_n7223_, new_n4717_, new_n8886_, new_n4718_,
    new_n8883_, new_n4719_, new_n8907_, new_n4720_, new_n8914_, new_n4721_,
    new_n8922_, new_n8789_, new_n4722_, new_n8926_, new_n4723_, new_n8936_,
    new_n4724_, new_n8948_, new_n4725_, new_n8945_, new_n4726_, new_n8963_,
    new_n7224_, new_n4727_, new_n8960_, new_n4728_, new_n8975_, new_n4729_,
    new_n8977_, new_n4730_, new_n8997_, new_n4731_, new_n9012_, new_n7225_,
    new_n4732_, new_n9009_, new_n4733_, new_n9019_, new_n4734_, new_n9023_,
    new_n4735_, new_n9033_, new_n4736_, new_n9039_, new_n7226_, new_n4737_,
    new_n9056_, new_n4738_, new_n9054_, new_n4739_, new_n9051_, new_n4740_,
    new_n9069_, new_n4741_, new_n9066_, new_n10704_, new_n9710_,
    new_n4742_, new_n9086_, new_n4743_, new_n9094_, new_n4744_, new_n9103_,
    new_n4745_, new_n9119_, new_n4746_, new_n9117_, new_n7227_, new_n4747_,
    new_n9114_, new_n4748_, new_n9132_, new_n4749_, new_n9129_, new_n4750_,
    new_n9140_, new_n4751_, new_n9149_, new_n7228_, new_n4752_, new_n9159_,
    new_n4753_, new_n9168_, new_n4754_, new_n9170_, new_n4755_, new_n9181_,
    new_n4756_, new_n9188_, new_n7229_, new_n4757_, new_n9193_, new_n4758_,
    new_n9204_, new_n4759_, new_n9211_, new_n4760_, new_n9213_, new_n4761_,
    new_n9224_, new_n7230_, new_n4762_, new_n9231_, new_n4763_, new_n9237_,
    new_n4764_, new_n9252_, new_n4765_, new_n9259_, new_n4766_, new_n9266_,
    new_n7231_, new_n4767_, new_n9286_, new_n4768_, new_n9308_, new_n4769_,
    new_n9317_, new_n4770_, new_n9324_, new_n4771_, new_n9332_, new_n7232_,
    new_n4772_, new_n9341_, new_n4773_, new_n9346_, new_n4774_, new_n9355_,
    new_n4775_, new_n9364_, new_n4776_, new_n9370_, new_n7233_, new_n4777_,
    new_n9379_, new_n4778_, new_n9385_, new_n4779_, new_n4780_, new_n9394_,
    new_n4781_, new_n9399_, new_n4782_, new_n7234_, new_n4783_, new_n9408_,
    new_n4784_, new_n9413_, new_n4785_, new_n9422_, new_n4786_, new_n9428_,
    new_n4787_, new_n9437_, new_n7235_, new_n4788_, new_n9443_, new_n4789_,
    new_n9452_, new_n4790_, new_n9458_, new_n4791_, new_n9467_, new_n4792_,
    new_n9473_, new_n7047_, new_n7236_, new_n4793_, new_n9481_, new_n4794_,
    new_n9488_, new_n4795_, new_n9497_, new_n4796_, new_n9502_, new_n4797_,
    new_n9511_, new_n7237_, new_n4798_, new_n9519_, new_n4799_, new_n9526_,
    new_n4800_, new_n9545_, new_n4801_, new_n9556_, new_n4802_, new_n9573_,
    new_n7238_, new_n4803_, new_n9577_, new_n4804_, new_n9587_, new_n4805_,
    new_n9591_, new_n4806_, new_n9602_, new_n4807_, new_n9606_, new_n7239_,
    new_n4808_, new_n9617_, new_n4809_, new_n9621_, new_n4810_, new_n9643_,
    new_n4811_, new_n9635_, new_n4812_, new_n9652_, new_n7240_, new_n4813_,
    new_n9656_, new_n4814_, new_n9667_, new_n4815_, new_n9678_, new_n4816_,
    new_n9682_, new_n4817_, new_n9690_, new_n7241_, new_n4818_, new_n9686_,
    new_n4819_, new_n9692_, new_n4820_, new_n9696_, new_n4821_, new_n9671_,
    new_n4822_, new_n9702_, new_n7242_, new_n4823_, new_n9706_, new_n4824_,
    new_n9715_, new_n4825_, new_n9719_, new_n4826_, new_n9731_, new_n4827_,
    new_n9743_, new_n7243_, new_n4828_, new_n9753_, new_n4829_, new_n9757_,
    new_n4830_, new_n9767_, new_n4831_, new_n9771_, new_n4832_, new_n9781_,
    new_n7244_, new_n4833_, new_n9785_, new_n4834_, new_n9795_, new_n4835_,
    new_n9799_, new_n4836_, new_n9808_, new_n4837_, new_n9820_, new_n7245_,
    new_n4838_, new_n9828_, new_n4839_, new_n9832_, new_n4840_, new_n9843_,
    new_n4841_, new_n9847_, new_n4842_, new_n9858_, new_n7048_, new_n7246_,
    new_n4843_, new_n9862_, new_n4844_, new_n9871_, new_n4845_, new_n9874_,
    new_n4846_, new_n9880_, new_n4847_, new_n9884_, new_n7247_, new_n4848_,
    new_n9891_, new_n4849_, new_n9908_, new_n4850_, new_n9895_, new_n4851_,
    new_n9917_, new_n4852_, new_n9921_, new_n7248_, new_n4853_, new_n9932_,
    new_n4854_, new_n9941_, new_n4855_, new_n9936_, new_n4856_, new_n9951_,
    new_n4857_, new_n9955_, new_n7249_, new_n4858_, new_n9962_, new_n4859_,
    new_n9966_, new_n4860_, new_n9977_, new_n4861_, new_n9981_, new_n4862_,
    new_n9991_, new_n7250_, new_n4863_, new_n10003_, new_n4864_,
    new_n10008_, new_n4865_, new_n10010_, new_n4866_, new_n10016_,
    new_n4867_, new_n10012_, new_n7251_, new_n4868_, new_n10018_,
    new_n4869_, new_n10024_, new_n4870_, new_n10020_, new_n4871_,
    new_n10026_, new_n4872_, new_n10036_, new_n7252_, new_n4873_,
    new_n10038_, new_n4874_, new_n10047_, new_n4875_, new_n10052_,
    new_n4876_, new_n10057_, new_n4877_, new_n10059_, new_n7253_,
    new_n4878_, new_n10072_, new_n4879_, new_n10074_, new_n4880_,
    new_n10051_, new_n4881_, new_n10077_, new_n4882_, new_n10079_,
    new_n7254_, new_n4883_, new_n10082_, new_n4884_, new_n10085_,
    new_n4885_, new_n10087_, new_n4886_, new_n10028_, new_n4887_,
    new_n10089_, new_n11129_, new_n4888_, new_n10092_, new_n4889_,
    new_n10098_, new_n4890_, new_n10100_, new_n4891_, new_n9995_,
    new_n4892_, new_n10105_, new_n7049_, new_n7255_, new_n4893_,
    new_n10112_, new_n4894_, new_n10133_, new_n4895_, new_n10131_,
    new_n4896_, new_n10141_, new_n4897_, new_n10143_, new_n9269_,
    new_n4898_, new_n10148_, new_n4899_, new_n10181_, new_n4900_,
    new_n10188_, new_n4901_, new_n10190_, new_n4902_, new_n10197_,
    new_n7256_, new_n4903_, new_n10203_, new_n4904_, new_n10205_,
    new_n4905_, new_n10211_, new_n4906_, new_n10213_, new_n4907_,
    new_n10216_, new_n7257_, new_n4908_, new_n10222_, new_n4909_,
    new_n10224_, new_n4910_, new_n10175_, new_n4911_, new_n10231_,
    new_n4912_, new_n10233_, new_n10135_, new_n4913_, new_n10236_,
    new_n4914_, new_n10238_, new_n4915_, new_n10244_, new_n4916_,
    new_n10246_, new_n4917_, new_n10249_, new_n7258_, new_n4918_,
    new_n10251_, new_n4919_, new_n10254_, new_n4920_, new_n10256_,
    new_n4921_, new_n10258_, new_n4922_, new_n10261_, new_n7259_,
    new_n4923_, new_n10264_, new_n4924_, new_n10266_, new_n4925_,
    new_n10269_, new_n4926_, new_n10272_, new_n4927_, new_n10274_,
    new_n10432_, new_n4928_, new_n10124_, new_n4929_, new_n10285_,
    new_n4930_, new_n10300_, new_n4931_, new_n10320_, new_n4932_,
    new_n10379_, new_n7260_, new_n4933_, new_n10392_, new_n4934_,
    new_n10400_, new_n4935_, new_n10386_, new_n4936_, new_n10330_,
    new_n4937_, new_n10428_, new_n7261_, new_n4938_, new_n10437_,
    new_n4939_, new_n10424_, new_n4940_, new_n10448_, new_n4941_,
    new_n10456_, new_n4942_, new_n10473_, new_n7050_, new_n7262_,
    new_n4943_, new_n10483_, new_n4944_, new_n10488_, new_n4945_,
    new_n10491_, new_n4946_, new_n10517_, new_n4947_, new_n10529_,
    new_n7263_, new_n4948_, new_n10555_, new_n4949_, new_n10575_,
    new_n4950_, new_n10579_, new_n4951_, new_n10588_, new_n4952_,
    new_n10591_, new_n7264_, new_n4953_, new_n10594_, new_n4954_,
    new_n10597_, new_n4955_, new_n10607_, new_n4956_, new_n10609_,
    new_n4957_, new_n10612_, new_n10316_, new_n4958_, new_n10615_,
    new_n4959_, new_n10618_, new_n4960_, new_n10534_, new_n4961_,
    new_n10622_, new_n4962_, new_n10639_, new_n7265_, new_n4963_,
    new_n10644_, new_n4964_, new_n10647_, new_n4965_, new_n10650_,
    new_n4966_, new_n10656_, new_n4967_, new_n10658_, new_n7266_,
    new_n4968_, new_n10661_, new_n4969_, new_n10665_, new_n4970_,
    new_n10669_, new_n4971_, new_n10671_, new_n4972_, new_n10673_,
    new_n7267_, new_n4973_, new_n10676_, new_n4974_, new_n10678_,
    new_n4975_, new_n10653_, new_n4976_, new_n10683_, new_n4977_,
    new_n10687_, new_n7268_, new_n4978_, new_n10690_, new_n4979_,
    new_n10692_, new_n4980_, new_n10695_, new_n4981_, new_n10710_,
    new_n4982_, new_n10719_, new_n7269_, new_n4983_, new_n10725_,
    new_n4984_, new_n10727_, new_n4985_, new_n10735_, new_n4986_,
    new_n10737_, new_n4987_, new_n10745_, new_n10323_, new_n4988_,
    new_n10747_, new_n4989_, new_n10753_, new_n4990_, new_n10755_,
    new_n4991_, new_n10766_, new_n4992_, new_n10768_, new_n7051_,
    new_n7270_, new_n4993_, new_n10774_, new_n4994_, new_n10776_,
    new_n4995_, new_n10787_, new_n4996_, new_n10789_, new_n4997_,
    new_n10795_, new_n8698_, new_n4998_, new_n10797_, new_n4999_,
    new_n10806_, new_n5000_, new_n10808_, new_n5001_, new_n10815_,
    new_n5002_, new_n10817_, new_n9625_, new_n5003_, new_n10827_,
    new_n5004_, new_n10829_, new_n5005_, new_n10835_, new_n5006_,
    new_n10837_, new_n5007_, new_n10848_, new_n7271_, new_n5008_,
    new_n10850_, new_n5009_, new_n10856_, new_n5010_, new_n10858_,
    new_n5011_, new_n10869_, new_n5012_, new_n10871_, new_n9484_,
    new_n5013_, new_n10877_, new_n5014_, new_n10879_, new_n5015_,
    new_n10889_, new_n5016_, new_n10891_, new_n5017_, new_n10897_,
    new_n7272_, new_n5018_, new_n10899_, new_n5019_, new_n10910_,
    new_n5020_, new_n10912_, new_n5021_, new_n10918_, new_n5022_,
    new_n10920_, new_n9790_, new_n5023_, new_n10931_, new_n5024_,
    new_n10933_, new_n5025_, new_n10939_, new_n5026_, new_n10941_,
    new_n5027_, new_n10952_, new_n7273_, new_n5028_, new_n10954_,
    new_n5029_, new_n10961_, new_n5030_, new_n10963_, new_n5031_,
    new_n10971_, new_n5032_, new_n10973_, new_n9903_, new_n5033_,
    new_n10979_, new_n5034_, new_n10981_, new_n5035_, new_n10988_,
    new_n5036_, new_n10990_, new_n5037_, new_n10996_, new_n7274_,
    new_n5038_, new_n10998_, new_n5039_, new_n11004_, new_n5040_,
    new_n11006_, new_n5041_, new_n11012_, new_n5042_, new_n11026_,
    new_n7052_, new_n9002_, new_n5043_, new_n11030_, new_n5044_,
    new_n11044_, new_n5045_, new_n11059_, new_n5046_, new_n11064_,
    new_n5047_, new_n11084_, new_n7275_, new_n5048_, new_n11112_,
    new_n5049_, new_n11118_, new_n5050_, new_n11124_, new_n5051_,
    new_n11127_, new_n5052_, new_n11128_, new_n11397_, new_n5053_,
    new_n11122_, new_n5054_, new_n11134_, new_n5055_, new_n11139_,
    new_n5056_, new_n11141_, new_n5057_, new_n11144_, new_n7276_,
    new_n5058_, new_n11147_, new_n5059_, new_n11150_, new_n5060_,
    new_n11100_, new_n5061_, new_n11157_, new_n5062_, new_n11177_,
    new_n9777_, new_n5063_, new_n11198_, new_n5064_, new_n11217_,
    new_n5065_, new_n11236_, new_n5066_, new_n11255_, new_n5067_,
    new_n11274_, new_n7277_, new_n5068_, new_n11295_, new_n5069_,
    new_n11305_, new_n5070_, new_n11311_, new_n5071_, new_n11314_,
    new_n5072_, new_n11317_, new_n9744_, new_n5073_, new_n11320_,
    new_n5074_, new_n11323_, new_n5075_, new_n11326_, new_n5076_,
    new_n11329_, new_n5077_, new_n11332_, new_n7278_, new_n5078_,
    new_n11335_, new_n5079_, new_n11338_, new_n5080_, new_n11342_,
    new_n5081_, new_n11350_, new_n5082_, new_n11354_, new_n9644_,
    new_n5083_, new_n11359_, new_n5084_, new_n11365_, new_n5085_,
    new_n11376_, new_n5086_, new_n11386_, new_n5087_, new_n11390_,
    new_n7279_, new_n5088_, new_n11394_, new_n5089_, new_n11402_,
    new_n5090_, new_n11412_, new_n5091_, new_n11418_, new_n5092_,
    new_n11422_, new_n9154_, new_n9561_, new_n5093_, new_n11425_,
    new_n5094_, new_n11429_, new_n5095_, new_n11438_, new_n5096_,
    new_n11443_, new_n5097_, new_n11448_, new_n7280_, new_n5098_,
    new_n11452_, new_n5099_, new_n11436_, new_n5100_, new_n11433_,
    new_n5101_, new_n11456_, new_n5102_, new_n11455_, new_n10465_,
    new_n5103_, new_n11462_, new_n5104_, new_n11466_, new_n5105_,
    new_n11469_, new_n5106_, new_n7573_, new_n5107_, new_n7575_,
    new_n7281_, new_n5108_, new_n7595_, new_n5109_, new_n7597_, new_n5110_,
    new_n7614_, new_n5111_, new_n7616_, new_n5112_, new_n7633_, new_n7282_,
    new_n5113_, new_n7635_, new_n5114_, new_n7648_, new_n5115_, new_n7654_,
    new_n5116_, new_n7656_, new_n5117_, new_n7676_, new_n11442_,
    new_n5118_, new_n7678_, new_n5119_, new_n7692_, new_n5120_, new_n7698_,
    new_n5121_, new_n7700_, new_n5122_, new_n7714_, new_n7283_, new_n5123_,
    new_n7717_, new_n5124_, new_n7720_, new_n5125_, new_n7723_, new_n5126_,
    new_n7726_, new_n5127_, new_n7727_, new_n10660_, new_n5128_,
    new_n7743_, new_n5129_, new_n7746_, new_n5130_, new_n7749_, new_n5131_,
    new_n7752_, new_n5132_, new_n7756_, new_n7284_, new_n5133_, new_n7760_,
    new_n5134_, new_n7764_, new_n5135_, new_n7771_, new_n5136_, new_n7779_,
    new_n5137_, new_n7787_, new_n10675_, new_n5138_, new_n7792_,
    new_n5139_, new_n7805_, new_n5140_, new_n7813_, new_n5141_, new_n7818_,
    new_n5142_, new_n7825_, new_n7053_, new_n7285_, new_n5143_, new_n7832_,
    new_n5144_, new_n7835_, new_n5145_, new_n7842_, new_n5146_, new_n7849_,
    new_n5147_, new_n7852_, new_n11352_, new_n5148_, new_n7859_,
    new_n5149_, new_n7866_, new_n5150_, new_n7869_, new_n5151_, new_n7876_,
    new_n5152_, new_n7883_, new_n7286_, new_n5153_, new_n7886_, new_n5154_,
    new_n7893_, new_n5155_, new_n7900_, new_n5156_, new_n7903_, new_n5157_,
    new_n7910_, new_n11368_, new_n5158_, new_n7917_, new_n5159_,
    new_n7920_, new_n5160_, new_n7927_, new_n5161_, new_n7934_, new_n5162_,
    new_n7937_, new_n7287_, new_n5163_, new_n7944_, new_n5164_, new_n7951_,
    new_n5165_, new_n7954_, new_n5166_, new_n7961_, new_n5167_, new_n7968_,
    new_n9241_, new_n5168_, new_n7971_, new_n5169_, new_n7978_, new_n5170_,
    new_n7985_, new_n5171_, new_n7988_, new_n5172_, new_n7995_, new_n7288_,
    new_n5173_, new_n8002_, new_n5174_, new_n8005_, new_n5175_, new_n8012_,
    new_n5176_, new_n8019_, new_n5177_, new_n8022_, new_n7289_, new_n5178_,
    new_n8029_, new_n5179_, new_n8036_, new_n5180_, new_n8039_, new_n5181_,
    new_n8046_, new_n5182_, new_n8053_, new_n9564_, new_n5183_, new_n8056_,
    new_n5184_, new_n8063_, new_n5185_, new_n8070_, new_n5186_, new_n8073_,
    new_n5187_, new_n8080_, new_n7290_, new_n5188_, new_n8087_, new_n5189_,
    new_n8090_, new_n5190_, new_n8097_, new_n5191_, new_n8104_, new_n5192_,
    new_n8107_, new_n7025_, new_n7054_, new_n7291_, new_n5193_, new_n8123_,
    new_n5194_, new_n8126_, new_n5195_, new_n8133_, new_n5196_, new_n8140_,
    new_n5197_, new_n8143_, new_n7292_, new_n5198_, new_n8158_, new_n5199_,
    new_n8161_, new_n5200_, new_n8168_, new_n5201_, new_n8175_, new_n5202_,
    new_n8178_, new_n7918_, new_n5203_, new_n8193_, new_n5204_, new_n8196_,
    new_n5205_, new_n8203_, new_n5206_, new_n8210_, new_n5207_, new_n8213_,
    new_n7293_, new_n5208_, new_n8227_, new_n5209_, new_n8229_, new_n5210_,
    new_n8236_, new_n5211_, new_n8243_, new_n5212_, new_n8246_, new_n7294_,
    new_n5213_, new_n8261_, new_n5214_, new_n8264_, new_n5215_, new_n8271_,
    new_n5216_, new_n8278_, new_n5217_, new_n8280_, new_n7295_, new_n5218_,
    new_n8285_, new_n5219_, new_n8294_, new_n5220_, new_n8298_, new_n5221_,
    new_n8403_, new_n5222_, new_n8411_, new_n11146_, new_n5223_,
    new_n8417_, new_n5224_, new_n8424_, new_n5225_, new_n8428_, new_n5226_,
    new_n8431_, new_n5227_, new_n8435_, new_n7296_, new_n5228_, new_n8448_,
    new_n5229_, new_n8453_, new_n5230_, new_n8461_, new_n5231_, new_n8463_,
    new_n5232_, new_n8469_, new_n9321_, new_n5233_, new_n8475_, new_n5234_,
    new_n8480_, new_n5235_, new_n8482_, new_n5236_, new_n8490_, new_n5237_,
    new_n8492_, new_n7297_, new_n5238_, new_n8500_, new_n5239_, new_n8505_,
    new_n5240_, new_n8510_, new_n5241_, new_n8526_, new_n5242_, new_n8528_,
    new_n10525_, new_n8517_, new_n5243_, new_n8534_, new_n5244_,
    new_n8538_, new_n5245_, new_n8543_, new_n5246_, new_n8550_, new_n5247_,
    new_n8558_, new_n7298_, new_n5248_, new_n8560_, new_n5249_, new_n8566_,
    new_n5250_, new_n8570_, new_n5251_, new_n8577_, new_n5252_, new_n8579_,
    new_n7299_, new_n5253_, new_n8588_, new_n5254_, new_n8593_, new_n5255_,
    new_n8595_, new_n5256_, new_n8603_, new_n5257_, new_n8605_, new_n7300_,
    new_n5258_, new_n8612_, new_n5259_, new_n8616_, new_n5260_, new_n8622_,
    new_n5261_, new_n8626_, new_n5262_, new_n8631_, new_n7301_, new_n5263_,
    new_n8636_, new_n5264_, new_n8644_, new_n5265_, new_n8646_, new_n5266_,
    new_n8651_, new_n5267_, new_n8654_, new_n7302_, new_n5268_, new_n8659_,
    new_n5269_, new_n8661_, new_n5270_, new_n8679_, new_n5271_, new_n8681_,
    new_n5272_, new_n8687_, new_n7303_, new_n5273_, new_n8703_, new_n5274_,
    new_n8705_, new_n5275_, new_n8712_, new_n5276_, new_n8716_, new_n5277_,
    new_n8721_, new_n7590_, new_n5278_, new_n8736_, new_n5279_, new_n8738_,
    new_n5280_, new_n8744_, new_n5281_, new_n8748_, new_n5282_, new_n8755_,
    new_n7304_, new_n5283_, new_n8757_, new_n5284_, new_n8764_, new_n5285_,
    new_n8769_, new_n5286_, new_n8771_, new_n5287_, new_n8782_, new_n7305_,
    new_n5288_, new_n8784_, new_n5289_, new_n8791_, new_n5290_, new_n8803_,
    new_n5291_, new_n8810_, new_n5292_, new_n8812_, new_n7055_, new_n7306_,
    new_n5293_, new_n8818_, new_n5294_, new_n8827_, new_n5295_, new_n8832_,
    new_n5296_, new_n8847_, new_n5297_, new_n8849_, new_n10436_,
    new_n5298_, new_n8855_, new_n5299_, new_n8859_, new_n5300_, new_n8864_,
    new_n5301_, new_n8866_, new_n5302_, new_n8874_, new_n7307_, new_n5303_,
    new_n8876_, new_n5304_, new_n8882_, new_n5305_, new_n8887_, new_n5306_,
    new_n8893_, new_n5307_, new_n8904_, new_n10686_, new_n5308_,
    new_n8906_, new_n5309_, new_n8913_, new_n5310_, new_n8925_, new_n5311_,
    new_n8933_, new_n5312_, new_n8935_, new_n7308_, new_n5313_, new_n8944_,
    new_n5314_, new_n8949_, new_n5315_, new_n8950_, new_n5316_, new_n8957_,
    new_n5317_, new_n8959_, new_n10664_, new_n5318_, new_n8965_,
    new_n5319_, new_n8974_, new_n5320_, new_n8978_, new_n5321_, new_n8994_,
    new_n5322_, new_n8996_, new_n7309_, new_n5323_, new_n8999_, new_n5324_,
    new_n9004_, new_n5325_, new_n9008_, new_n5326_, new_n9013_, new_n5327_,
    new_n9022_, new_n8624_, new_n5328_, new_n9030_, new_n5329_, new_n9032_,
    new_n5330_, new_n9038_, new_n5331_, new_n9041_, new_n5332_, new_n9048_,
    new_n7310_, new_n5333_, new_n9050_, new_n5334_, new_n9065_, new_n5335_,
    new_n9070_, new_n5336_, new_n9072_, new_n5337_, new_n9083_, new_n7311_,
    new_n5338_, new_n9085_, new_n5339_, new_n9093_, new_n5340_, new_n9104_,
    new_n5341_, new_n9105_, new_n5342_, new_n9111_, new_n7056_, new_n7312_,
    new_n5343_, new_n9113_, new_n5344_, new_n9128_, new_n5345_, new_n9134_,
    new_n5346_, new_n9146_, new_n5347_, new_n9148_, new_n11461_,
    new_n5348_, new_n9151_, new_n5349_, new_n9158_, new_n5350_, new_n9169_,
    new_n5351_, new_n9178_, new_n5352_, new_n9180_, new_n7313_, new_n5353_,
    new_n9187_, new_n5354_, new_n9194_, new_n5355_, new_n9201_, new_n5356_,
    new_n9203_, new_n5357_, new_n9210_, new_n7314_, new_n5358_, new_n9214_,
    new_n5359_, new_n9221_, new_n5360_, new_n9223_, new_n5361_, new_n9230_,
    new_n5362_, new_n9236_, new_n7315_, new_n5363_, new_n9249_, new_n5364_,
    new_n9251_, new_n5365_, new_n9258_, new_n5366_, new_n9264_, new_n5367_,
    new_n9268_, new_n7316_, new_n5368_, new_n9273_, new_n5369_, new_n9277_,
    new_n5370_, new_n9310_, new_n5371_, new_n9326_, new_n5372_, new_n9334_,
    new_n7317_, new_n5373_, new_n9348_, new_n5374_, new_n9357_, new_n5375_,
    new_n9372_, new_n5376_, new_n9387_, new_n5377_, new_n9401_, new_n7318_,
    new_n5378_, new_n9415_, new_n5379_, new_n9430_, new_n5380_, new_n9445_,
    new_n5381_, new_n9460_, new_n5382_, new_n9475_, new_n7319_, new_n5383_,
    new_n9490_, new_n5384_, new_n9504_, new_n5385_, new_n9513_, new_n5386_,
    new_n9528_, new_n5387_, new_n9546_, new_n7320_, new_n5388_, new_n9550_,
    new_n5389_, new_n9557_, new_n5390_, new_n9572_, new_n5391_, new_n9574_,
    new_n5392_, new_n9576_, new_n7608_, new_n7321_, new_n5393_, new_n9588_,
    new_n5394_, new_n9590_, new_n5395_, new_n9601_, new_n5396_, new_n9603_,
    new_n5397_, new_n9605_, new_n7322_, new_n5398_, new_n9618_, new_n5399_,
    new_n9620_, new_n5400_, new_n9630_, new_n5401_, new_n9634_, new_n5402_,
    new_n9653_, new_n7323_, new_n5403_, new_n9655_, new_n5404_, new_n9666_,
    new_n5405_, new_n9668_, new_n5406_, new_n9670_, new_n5407_, new_n9679_,
    new_n7324_, new_n5408_, new_n9683_, new_n5409_, new_n9687_, new_n5410_,
    new_n9691_, new_n5411_, new_n9703_, new_n5412_, new_n9705_, new_n7325_,
    new_n5413_, new_n9716_, new_n5414_, new_n9718_, new_n5415_, new_n9730_,
    new_n5416_, new_n9732_, new_n5417_, new_n9734_, new_n7326_, new_n5418_,
    new_n9739_, new_n5419_, new_n9754_, new_n5420_, new_n9756_, new_n5421_,
    new_n9766_, new_n5422_, new_n9768_, new_n7327_, new_n5423_, new_n9770_,
    new_n5424_, new_n9782_, new_n5425_, new_n9784_, new_n5426_, new_n9796_,
    new_n5427_, new_n9798_, new_n7328_, new_n5428_, new_n9809_, new_n5429_,
    new_n9811_, new_n5430_, new_n9816_, new_n5431_, new_n9827_, new_n5432_,
    new_n9829_, new_n7329_, new_n5433_, new_n9831_, new_n5434_, new_n9844_,
    new_n5435_, new_n9846_, new_n5436_, new_n9859_, new_n5437_, new_n9861_,
    new_n7330_, new_n5438_, new_n9872_, new_n5439_, new_n9875_, new_n5440_,
    new_n9879_, new_n5441_, new_n9881_, new_n5442_, new_n9883_, new_n7057_,
    new_n7331_, new_n5443_, new_n9892_, new_n5444_, new_n9894_, new_n5445_,
    new_n9901_, new_n5446_, new_n9910_, new_n5447_, new_n9916_, new_n7332_,
    new_n5448_, new_n9918_, new_n5449_, new_n9920_, new_n5450_, new_n9933_,
    new_n5451_, new_n9935_, new_n5452_, new_n9938_, new_n7333_, new_n5453_,
    new_n9947_, new_n5454_, new_n9952_, new_n5455_, new_n9954_, new_n5456_,
    new_n9963_, new_n5457_, new_n9965_, new_n8800_, new_n5458_, new_n9978_,
    new_n5459_, new_n9980_, new_n5460_, new_n9985_, new_n5461_, new_n9990_,
    new_n5462_, new_n9992_, new_n7334_, new_n5463_, new_n9994_, new_n5464_,
    new_n10009_, new_n5465_, new_n10011_, new_n5466_, new_n10013_,
    new_n5467_, new_n10017_, new_n9101_, new_n5468_, new_n10019_,
    new_n5469_, new_n10021_, new_n5470_, new_n10025_, new_n5471_,
    new_n10027_, new_n5472_, new_n10029_, new_n7335_, new_n5473_,
    new_n10037_, new_n5474_, new_n10039_, new_n5475_, new_n10045_,
    new_n5476_, new_n10058_, new_n5477_, new_n10060_, new_n7336_,
    new_n5478_, new_n10066_, new_n5479_, new_n10073_, new_n5480_,
    new_n10075_, new_n5481_, new_n10078_, new_n5482_, new_n10080_,
    new_n7337_, new_n5483_, new_n10083_, new_n5484_, new_n10086_,
    new_n5485_, new_n10088_, new_n5486_, new_n10090_, new_n5487_,
    new_n10093_, new_n7338_, new_n5488_, new_n10099_, new_n5489_,
    new_n10101_, new_n5490_, new_n10106_, new_n5491_, new_n10111_,
    new_n5492_, new_n10113_, new_n8892_, new_n10740_, new_n5493_,
    new_n10120_, new_n5494_, new_n10129_, new_n5495_, new_n10142_,
    new_n5496_, new_n10144_, new_n5497_, new_n10146_, new_n10761_,
    new_n5498_, new_n10160_, new_n5499_, new_n10167_, new_n5500_,
    new_n10179_, new_n5501_, new_n10189_, new_n5502_, new_n10191_,
    new_n7339_, new_n5503_, new_n10193_, new_n5504_, new_n10198_,
    new_n5505_, new_n10204_, new_n5506_, new_n10206_, new_n5507_,
    new_n10212_, new_n10843_, new_n5508_, new_n10214_, new_n5509_,
    new_n10217_, new_n5510_, new_n10223_, new_n5511_, new_n10225_,
    new_n5512_, new_n10232_, new_n7340_, new_n5513_, new_n10234_,
    new_n5514_, new_n10237_, new_n5515_, new_n10239_, new_n5516_,
    new_n10245_, new_n5517_, new_n10247_, new_n10905_, new_n5518_,
    new_n10250_, new_n5519_, new_n10252_, new_n5520_, new_n10255_,
    new_n5521_, new_n10257_, new_n5522_, new_n10259_, new_n7341_,
    new_n5523_, new_n10262_, new_n5524_, new_n10265_, new_n5525_,
    new_n10267_, new_n5526_, new_n5527_, new_n10270_, new_n5528_,
    new_n10926_, new_n10273_, new_n5529_, new_n10275_, new_n5530_,
    new_n10276_, new_n5531_, new_n10280_, new_n5532_, new_n10286_,
    new_n5533_, new_n7342_, new_n10301_, new_n5534_, new_n10335_,
    new_n5535_, new_n10339_, new_n5536_, new_n10373_, new_n5537_,
    new_n10387_, new_n5538_, new_n7343_, new_n10408_, new_n5539_,
    new_n10425_, new_n5540_, new_n10429_, new_n5541_, new_n10438_,
    new_n5542_, new_n10449_, new_n5543_, new_n7058_, new_n10966_,
    new_n10457_, new_n5544_, new_n10469_, new_n5545_, new_n10474_,
    new_n5546_, new_n10477_, new_n5547_, new_n10481_, new_n5548_,
    new_n7344_, new_n10490_, new_n5549_, new_n10492_, new_n5550_,
    new_n10494_, new_n5551_, new_n10499_, new_n5552_, new_n10500_,
    new_n5553_, new_n7345_, new_n10502_, new_n5554_, new_n10505_,
    new_n5555_, new_n10508_, new_n5556_, new_n10513_, new_n5557_,
    new_n10524_, new_n5558_, new_n7346_, new_n10526_, new_n5559_,
    new_n10528_, new_n5560_, new_n10530_, new_n5561_, new_n10535_,
    new_n5562_, new_n10543_, new_n5563_, new_n8685_, new_n10550_,
    new_n5564_, new_n10552_, new_n5565_, new_n10559_, new_n5566_,
    new_n10567_, new_n5567_, new_n10570_, new_n5568_, new_n7347_,
    new_n10573_, new_n5569_, new_n10574_, new_n5570_, new_n10585_,
    new_n5571_, new_n10623_, new_n5572_, new_n10627_, new_n5573_,
    new_n7348_, new_n10629_, new_n5574_, new_n10631_, new_n5575_,
    new_n10642_, new_n5576_, new_n10654_, new_n5577_, new_n10708_,
    new_n5578_, new_n7349_, new_n10718_, new_n5579_, new_n10726_,
    new_n5580_, new_n10728_, new_n5581_, new_n10736_, new_n5582_,
    new_n10738_, new_n5583_, new_n7350_, new_n10746_, new_n5584_,
    new_n10748_, new_n5585_, new_n10754_, new_n5586_, new_n10756_,
    new_n5587_, new_n10760_, new_n5588_, new_n7783_, new_n10767_,
    new_n5589_, new_n10769_, new_n5590_, new_n10775_, new_n5591_,
    new_n10777_, new_n5592_, new_n10782_, new_n5593_, new_n7059_,
    new_n7351_, new_n10788_, new_n5594_, new_n10790_, new_n5595_,
    new_n10796_, new_n5596_, new_n10798_, new_n5597_, new_n10807_,
    new_n5598_, new_n7352_, new_n10809_, new_n5599_, new_n10816_,
    new_n5600_, new_n10818_, new_n5601_, new_n5602_, new_n10828_,
    new_n5603_, new_n10830_, new_n8439_, new_n5604_, new_n10836_,
    new_n5605_, new_n10838_, new_n5606_, new_n10842_, new_n5607_,
    new_n10849_, new_n5608_, new_n10851_, new_n7353_, new_n5609_,
    new_n10857_, new_n5610_, new_n10859_, new_n5611_, new_n10864_,
    new_n5612_, new_n10870_, new_n5613_, new_n10872_, new_n7354_,
    new_n5614_, new_n10878_, new_n5615_, new_n10880_, new_n5616_,
    new_n10890_, new_n5617_, new_n10892_, new_n5618_, new_n10898_,
    new_n7355_, new_n5619_, new_n10900_, new_n5620_, new_n10904_,
    new_n5621_, new_n10911_, new_n5622_, new_n10913_, new_n5623_,
    new_n10919_, new_n10822_, new_n5624_, new_n10921_, new_n5625_,
    new_n10925_, new_n5626_, new_n10932_, new_n5627_, new_n10934_,
    new_n5628_, new_n10940_, new_n7356_, new_n5629_, new_n10942_,
    new_n5630_, new_n10947_, new_n5631_, new_n10953_, new_n5632_,
    new_n10955_, new_n5633_, new_n10962_, new_n7357_, new_n5634_,
    new_n10964_, new_n5635_, new_n10972_, new_n5636_, new_n10974_,
    new_n5637_, new_n10980_, new_n5638_, new_n10982_, new_n7358_,
    new_n5639_, new_n10989_, new_n5640_, new_n10991_, new_n5641_,
    new_n10997_, new_n5642_, new_n10999_, new_n5643_, new_n11005_,
    new_n11269_, new_n7359_, new_n5644_, new_n11007_, new_n5645_,
    new_n11013_, new_n5646_, new_n11027_, new_n5647_, new_n11043_,
    new_n5648_, new_n11045_, new_n7360_, new_n5649_, new_n11063_,
    new_n5650_, new_n11065_, new_n5651_, new_n11085_, new_n5652_,
    new_n11097_, new_n5653_, new_n11101_, new_n7361_, new_n5654_,
    new_n11111_, new_n5655_, new_n11121_, new_n5656_, new_n11125_,
    new_n5657_, new_n11131_, new_n5658_, new_n11135_, new_n7362_,
    new_n5659_, new_n11140_, new_n5660_, new_n11142_, new_n5661_,
    new_n11156_, new_n5662_, new_n11158_, new_n5663_, new_n11176_,
    new_n7363_, new_n5664_, new_n11178_, new_n5665_, new_n11191_,
    new_n5666_, new_n11197_, new_n5667_, new_n11199_, new_n5668_,
    new_n11216_, new_n11033_, new_n5669_, new_n11218_, new_n5670_,
    new_n11235_, new_n5671_, new_n11237_, new_n5672_, new_n11254_,
    new_n5673_, new_n11256_, new_n7364_, new_n5674_, new_n11273_,
    new_n5675_, new_n11275_, new_n5676_, new_n11293_, new_n5677_,
    new_n11296_, new_n5678_, new_n11309_, new_n7365_, new_n5679_,
    new_n11312_, new_n5680_, new_n11315_, new_n5681_, new_n11318_,
    new_n5682_, new_n11321_, new_n5683_, new_n11324_, new_n7366_,
    new_n5684_, new_n11327_, new_n5685_, new_n11330_, new_n5686_,
    new_n11333_, new_n5687_, new_n11336_, new_n5688_, new_n11339_,
    new_n7367_, new_n5689_, new_n11343_, new_n5690_, new_n11348_,
    new_n5691_, new_n11353_, new_n5692_, new_n11369_, new_n5693_,
    new_n11380_, new_n7026_, new_n7060_, new_n7368_, new_n5694_,
    new_n11383_, new_n5695_, new_n11387_, new_n5696_, new_n11389_,
    new_n5697_, new_n11395_, new_n5698_, new_n11405_, new_n7369_,
    new_n5699_, new_n11413_, new_n5700_, new_n11416_, new_n5701_,
    new_n11419_, new_n5702_, new_n11423_, new_n5703_, new_n11426_,
    new_n7370_, new_n5704_, new_n11430_, new_n5705_, new_n11470_,
    new_n5706_, new_n7577_, new_n5707_, new_n7583_, new_n5708_, new_n7598_,
    new_n7371_, new_n5709_, new_n7618_, new_n5710_, new_n7623_, new_n5711_,
    new_n7636_, new_n5712_, new_n7638_, new_n5713_, new_n7658_, new_n7372_,
    new_n5714_, new_n7660_, new_n5715_, new_n7665_, new_n5716_, new_n7667_,
    new_n5717_, new_n7679_, new_n5718_, new_n7681_, new_n7373_, new_n5719_,
    new_n7702_, new_n5720_, new_n7704_, new_n5721_, new_n7709_, new_n5722_,
    new_n7711_, new_n5723_, new_n7801_, new_n7374_, new_n5724_, new_n7821_,
    new_n5725_, new_n7838_, new_n5726_, new_n7855_, new_n5727_, new_n7872_,
    new_n5728_, new_n7889_, new_n7375_, new_n5729_, new_n7906_, new_n5730_,
    new_n7923_, new_n5731_, new_n7940_, new_n5732_, new_n7957_, new_n5733_,
    new_n7974_, new_n7376_, new_n5734_, new_n7991_, new_n5735_, new_n8008_,
    new_n5736_, new_n8025_, new_n5737_, new_n8042_, new_n5738_, new_n8059_,
    new_n7377_, new_n5739_, new_n8076_, new_n5740_, new_n8093_, new_n5741_,
    new_n8110_, new_n5742_, new_n8129_, new_n5743_, new_n8146_,
    new_n11172_, new_n7378_, new_n5744_, new_n8164_, new_n5745_,
    new_n8181_, new_n5746_, new_n8199_, new_n5747_, new_n8216_, new_n5748_,
    new_n8232_, new_n7379_, new_n5749_, new_n8249_, new_n5750_, new_n8267_,
    new_n5751_, new_n8302_, new_n5752_, new_n8306_, new_n5753_, new_n8309_,
    new_n7380_, new_n5754_, new_n8312_, new_n5755_, new_n8315_, new_n5756_,
    new_n8318_, new_n5757_, new_n8321_, new_n5758_, new_n8324_, new_n7381_,
    new_n5759_, new_n8327_, new_n5760_, new_n8330_, new_n5761_, new_n8333_,
    new_n5762_, new_n8336_, new_n5763_, new_n8339_, new_n7382_, new_n5764_,
    new_n8342_, new_n5765_, new_n8345_, new_n5766_, new_n8348_, new_n5767_,
    new_n8351_, new_n5768_, new_n8354_, new_n7383_, new_n5769_, new_n8357_,
    new_n5770_, new_n8360_, new_n5771_, new_n8363_, new_n5772_, new_n8366_,
    new_n5773_, new_n8369_, new_n7384_, new_n5774_, new_n8372_, new_n5775_,
    new_n8375_, new_n5776_, new_n8378_, new_n5777_, new_n8381_, new_n5778_,
    new_n8384_, new_n7947_, new_n5779_, new_n8387_, new_n5780_, new_n8390_,
    new_n5781_, new_n8393_, new_n5782_, new_n8396_, new_n5783_, new_n8401_,
    new_n7385_, new_n5784_, new_n8409_, new_n5785_, new_n8421_, new_n5786_,
    new_n8458_, new_n5787_, new_n8484_, new_n5788_, new_n8487_, new_n7386_,
    new_n5789_, new_n8523_, new_n5790_, new_n8555_, new_n5791_, new_n8574_,
    new_n5792_, new_n8600_, new_n5793_, new_n8638_, new_n7061_, new_n7387_,
    new_n5794_, new_n8641_, new_n5795_, new_n8676_, new_n5796_, new_n8700_,
    new_n5797_, new_n8733_, new_n5798_, new_n8749_, new_n10410_,
    new_n5799_, new_n8752_, new_n5800_, new_n8773_, new_n5801_, new_n8779_,
    new_n5802_, new_n8807_, new_n5803_, new_n8844_, new_n7388_, new_n5804_,
    new_n8868_, new_n5805_, new_n8871_, new_n5806_, new_n8901_, new_n5807_,
    new_n8930_, new_n5808_, new_n8951_, new_n10338_, new_n5809_,
    new_n8954_, new_n5810_, new_n8983_, new_n5811_, new_n8991_, new_n5812_,
    new_n9027_, new_n5813_, new_n9042_, new_n7389_, new_n5814_, new_n9045_,
    new_n5815_, new_n9062_, new_n5816_, new_n9074_, new_n5817_, new_n9080_,
    new_n5818_, new_n9108_, new_n7390_, new_n5819_, new_n9123_, new_n5820_,
    new_n9143_, new_n5821_, new_n9175_, new_n5822_, new_n9198_, new_n5823_,
    new_n9215_, new_n7391_, new_n5824_, new_n9218_, new_n5825_, new_n9246_,
    new_n5826_, new_n9262_, new_n5827_, new_n9289_, new_n5828_, new_n9291_,
    new_n7392_, new_n5829_, new_n9295_, new_n5830_, new_n9298_, new_n5831_,
    new_n9307_, new_n5832_, new_n9316_, new_n5833_, new_n9323_,
    new_n10445_, new_n5834_, new_n9327_, new_n5835_, new_n9331_,
    new_n5836_, new_n9335_, new_n5837_, new_n9340_, new_n5838_, new_n9345_,
    new_n7393_, new_n5839_, new_n9349_, new_n5840_, new_n9354_, new_n5841_,
    new_n9358_, new_n5842_, new_n9363_, new_n5843_, new_n9369_, new_n7062_,
    new_n7394_, new_n5844_, new_n9373_, new_n5845_, new_n9378_, new_n5846_,
    new_n9384_, new_n5847_, new_n9388_, new_n5848_, new_n9393_, new_n7913_,
    new_n5849_, new_n9398_, new_n5850_, new_n9402_, new_n5851_, new_n9407_,
    new_n5852_, new_n9412_, new_n5853_, new_n9416_, new_n7395_, new_n5854_,
    new_n9421_, new_n5855_, new_n9427_, new_n5856_, new_n9431_, new_n5857_,
    new_n9436_, new_n5858_, new_n9442_, new_n7396_, new_n5859_, new_n9446_,
    new_n5860_, new_n9451_, new_n5861_, new_n9457_, new_n5862_, new_n9461_,
    new_n5863_, new_n9466_, new_n7397_, new_n5864_, new_n9472_, new_n5865_,
    new_n9476_, new_n5866_, new_n9480_, new_n5867_, new_n9487_, new_n5868_,
    new_n9491_, new_n7398_, new_n5869_, new_n9496_, new_n5870_, new_n9501_,
    new_n5871_, new_n9505_, new_n5872_, new_n9510_, new_n5873_, new_n9514_,
    new_n7399_, new_n5874_, new_n9518_, new_n5875_, new_n9525_, new_n5876_,
    new_n9529_, new_n5877_, new_n9534_, new_n5878_, new_n9535_, new_n7400_,
    new_n5879_, new_n9559_, new_n5880_, new_n10046_, new_n5881_,
    new_n10153_, new_n5882_, new_n10161_, new_n5883_, new_n10162_,
    new_n7401_, new_n5884_, new_n10168_, new_n5885_, new_n10180_,
    new_n5886_, new_n10226_, new_n5887_, new_n10287_, new_n5888_,
    new_n10289_, new_n9352_, new_n5889_, new_n10293_, new_n5890_,
    new_n10295_, new_n5891_, new_n10302_, new_n5892_, new_n10304_,
    new_n5893_, new_n10309_, new_n9823_, new_n7402_, new_n5894_,
    new_n10311_, new_n5895_, new_n10326_, new_n5896_, new_n10327_,
    new_n5897_, new_n10341_, new_n5898_, new_n10343_, new_n7403_,
    new_n5899_, new_n10345_, new_n5900_, new_n10347_, new_n5901_,
    new_n10349_, new_n5902_, new_n10351_, new_n5903_, new_n10353_,
    new_n9522_, new_n5904_, new_n10354_, new_n5905_, new_n10356_,
    new_n5906_, new_n10358_, new_n5907_, new_n10360_, new_n5908_,
    new_n10362_, new_n7404_, new_n5909_, new_n10364_, new_n5910_,
    new_n10366_, new_n5911_, new_n10368_, new_n5912_, new_n10394_,
    new_n5913_, new_n10475_, new_n9761_, new_n5914_, new_n10476_,
    new_n5915_, new_n10485_, new_n5916_, new_n10532_, new_n5917_,
    new_n10533_, new_n5918_, new_n10545_, new_n7405_, new_n5919_,
    new_n10547_, new_n5920_, new_n10548_, new_n5921_, new_n10557_,
    new_n5922_, new_n10560_, new_n5923_, new_n10571_, new_n7406_,
    new_n5924_, new_n10576_, new_n5925_, new_n10577_, new_n5926_,
    new_n10581_, new_n5927_, new_n10624_, new_n5928_, new_n10645_,
    new_n8416_, new_n5929_, new_n10646_, new_n5930_, new_n5931_,
    new_n5932_, new_n10706_, new_n5933_, new_n10716_, new_n5934_,
    new_n10722_, new_n7407_, new_n5935_, new_n10732_, new_n5936_,
    new_n10742_, new_n5937_, new_n10750_, new_n5938_, new_n10763_,
    new_n5939_, new_n10771_, new_n7408_, new_n5940_, new_n10784_,
    new_n5941_, new_n10792_, new_n5942_, new_n10803_, new_n5943_,
    new_n10812_, new_n5944_, new_n10824_, new_n7063_, new_n7409_,
    new_n5945_, new_n10832_, new_n5946_, new_n10845_, new_n5947_,
    new_n10853_, new_n5948_, new_n10866_, new_n5949_, new_n10874_,
    new_n7410_, new_n5950_, new_n10886_, new_n5951_, new_n10894_,
    new_n5952_, new_n10907_, new_n5953_, new_n10915_, new_n5954_,
    new_n10928_, new_n7411_, new_n5955_, new_n10936_, new_n5956_,
    new_n10949_, new_n5957_, new_n10958_, new_n5958_, new_n10968_,
    new_n5959_, new_n10976_, new_n7412_, new_n5960_, new_n10985_,
    new_n5961_, new_n10993_, new_n5962_, new_n11001_, new_n5963_,
    new_n11009_, new_n5964_, new_n11046_, new_n10419_, new_n5965_,
    new_n11048_, new_n5966_, new_n11053_, new_n5967_, new_n11055_,
    new_n5968_, new_n11067_, new_n5969_, new_n11069_, new_n7413_,
    new_n5970_, new_n11086_, new_n5971_, new_n11088_, new_n5972_,
    new_n11160_, new_n5973_, new_n11162_, new_n5974_, new_n11168_,
    new_n7414_, new_n5975_, new_n11180_, new_n5976_, new_n11182_,
    new_n5977_, new_n11200_, new_n5978_, new_n11202_, new_n5979_,
    new_n11207_, new_n10409_, new_n5980_, new_n11209_, new_n5981_,
    new_n11219_, new_n5982_, new_n11221_, new_n5983_, new_n11238_,
    new_n5984_, new_n11240_, new_n7415_, new_n5985_, new_n11244_,
    new_n5986_, new_n11246_, new_n5987_, new_n11257_, new_n5988_,
    new_n11259_, new_n5989_, new_n11276_, new_n7416_, new_n5990_,
    new_n11278_, new_n5991_, new_n11284_, new_n5992_, new_n11286_,
    new_n5993_, new_n11297_, new_n5994_, new_n11299_, new_n9693_,
    new_n7417_, new_n5995_, new_n5996_, new_n11367_, new_n5997_,
    new_n5998_, new_n5999_, new_n11440_, new_n6000_, new_n11458_,
    new_n6001_, new_n7418_, new_n7578_, new_n6002_, new_n7604_, new_n6003_,
    new_n7606_, new_n6004_, new_n7619_, new_n6005_, new_n6006_, new_n7647_,
    new_n8776_, new_n6007_, new_n7659_, new_n6008_, new_n6009_, new_n7691_,
    new_n6010_, new_n7703_, new_n6011_, new_n7721_, new_n6012_, new_n7419_,
    new_n7800_, new_n6013_, new_n7820_, new_n6014_, new_n7837_, new_n6015_,
    new_n7854_, new_n6016_, new_n7871_, new_n6017_, new_n9077_, new_n7888_,
    new_n6018_, new_n7905_, new_n6019_, new_n7922_, new_n6020_, new_n7939_,
    new_n6021_, new_n7956_, new_n6022_, new_n7420_, new_n7973_, new_n6023_,
    new_n7990_, new_n6024_, new_n8007_, new_n6025_, new_n8024_, new_n6026_,
    new_n8041_, new_n6027_, new_n9141_, new_n8058_, new_n6028_, new_n8075_,
    new_n6029_, new_n8092_, new_n6030_, new_n8109_, new_n6031_, new_n8128_,
    new_n6032_, new_n7421_, new_n8145_, new_n6033_, new_n8163_, new_n6034_,
    new_n8180_, new_n6035_, new_n8198_, new_n6036_, new_n8215_, new_n6037_,
    new_n10418_, new_n8231_, new_n6038_, new_n8248_, new_n6039_,
    new_n8266_, new_n6040_, new_n8301_, new_n6041_, new_n8305_, new_n6042_,
    new_n7422_, new_n8308_, new_n6043_, new_n8311_, new_n6044_, new_n8314_,
    new_n6045_, new_n8317_, new_n6046_, new_n8320_, new_n6047_, new_n7064_,
    new_n7423_, new_n8323_, new_n6048_, new_n8326_, new_n6049_, new_n8329_,
    new_n6050_, new_n8332_, new_n6051_, new_n8335_, new_n6052_, new_n7424_,
    new_n8338_, new_n6053_, new_n8341_, new_n6054_, new_n8344_, new_n6055_,
    new_n8347_, new_n6056_, new_n8350_, new_n6057_, new_n9185_, new_n8353_,
    new_n6058_, new_n8356_, new_n6059_, new_n8359_, new_n6060_, new_n8362_,
    new_n6061_, new_n8365_, new_n6062_, new_n7425_, new_n8368_, new_n6063_,
    new_n8371_, new_n6064_, new_n8374_, new_n6065_, new_n8377_, new_n6066_,
    new_n8380_, new_n6067_, new_n7426_, new_n8383_, new_n6068_, new_n8386_,
    new_n6069_, new_n8389_, new_n6070_, new_n8392_, new_n6071_, new_n8395_,
    new_n6072_, new_n7427_, new_n8400_, new_n6073_, new_n8408_, new_n6074_,
    new_n8436_, new_n6075_, new_n8420_, new_n6076_, new_n8457_, new_n6077_,
    new_n7428_, new_n8514_, new_n6078_, new_n8486_, new_n6079_, new_n8522_,
    new_n6080_, new_n8571_, new_n6081_, new_n8554_, new_n6082_, new_n7429_,
    new_n8573_, new_n6083_, new_n6084_, new_n8599_, new_n6085_, new_n8640_,
    new_n6086_, new_n6087_, new_n8675_, new_n6088_, new_n7430_, new_n8699_,
    new_n6089_, new_n8732_, new_n6090_, new_n8772_, new_n6091_, new_n8751_,
    new_n6092_, new_n8778_, new_n6093_, new_n10882_, new_n8819_,
    new_n6094_, new_n8823_, new_n6095_, new_n8825_, new_n6096_, new_n8842_,
    new_n6097_, new_n8806_, new_n6098_, new_n9244_, new_n8404_, new_n8843_,
    new_n6099_, new_n8870_, new_n6100_, new_n8900_, new_n6101_, new_n8929_,
    new_n6102_, new_n8966_, new_n6103_, new_n7431_, new_n8970_, new_n6104_,
    new_n8953_, new_n6105_, new_n9000_, new_n6106_, new_n8990_, new_n6107_,
    new_n9026_, new_n6108_, new_n11022_, new_n9058_, new_n6109_,
    new_n9073_, new_n6110_, new_n9044_, new_n6111_, new_n9079_, new_n6112_,
    new_n9124_, new_n6113_, new_n7432_, new_n9107_, new_n6114_, new_n9152_,
    new_n6115_, new_n9142_, new_n6116_, new_n9174_, new_n6117_, new_n9197_,
    new_n6118_, new_n7433_, new_n9217_, new_n6119_, new_n9245_, new_n6120_,
    new_n9270_, new_n6121_, new_n9271_, new_n6122_, new_n9261_, new_n6123_,
    new_n7434_, new_n9288_, new_n6124_, new_n9294_, new_n6125_, new_n9297_,
    new_n6126_, new_n9301_, new_n6127_, new_n9328_, new_n6128_, new_n7435_,
    new_n9337_, new_n6129_, new_n9360_, new_n6130_, new_n9375_, new_n6131_,
    new_n9390_, new_n6132_, new_n9404_, new_n6133_, new_n7436_, new_n9418_,
    new_n6134_, new_n9433_, new_n6135_, new_n9448_, new_n6136_, new_n9463_,
    new_n6137_, new_n9477_, new_n6138_, new_n7437_, new_n9493_, new_n6139_,
    new_n9507_, new_n6140_, new_n9515_, new_n6141_, new_n9531_, new_n6142_,
    new_n9533_, new_n6143_, new_n7438_, new_n10067_, new_n6144_,
    new_n10136_, new_n6145_, new_n6146_, new_n10147_, new_n6147_,
    new_n10288_, new_n6148_, new_n10294_, new_n7065_, new_n7439_,
    new_n6149_, new_n10303_, new_n6150_, new_n10310_, new_n6151_,
    new_n6152_, new_n10380_, new_n6153_, new_n10395_, new_n6154_,
    new_n7440_, new_n6155_, new_n10328_, new_n6156_, new_n6157_,
    new_n10480_, new_n6158_, new_n10484_, new_n6159_, new_n6160_,
    new_n6161_, new_n7441_, new_n6162_, new_n6163_, new_n6164_,
    new_n10580_, new_n6165_, new_n6166_, new_n6167_, new_n6168_,
    new_n10689_, new_n6169_, new_n7442_, new_n10325_, new_n6170_,
    new_n10705_, new_n6171_, new_n10715_, new_n6172_, new_n10721_,
    new_n6173_, new_n10731_, new_n6174_, new_n7443_, new_n10741_,
    new_n6175_, new_n10749_, new_n6176_, new_n10762_, new_n6177_,
    new_n10770_, new_n6178_, new_n10783_, new_n6179_, new_n9290_,
    new_n10791_, new_n6180_, new_n10802_, new_n6181_, new_n10811_,
    new_n6182_, new_n10823_, new_n6183_, new_n10831_, new_n6184_,
    new_n7444_, new_n10844_, new_n6185_, new_n10852_, new_n6186_,
    new_n10865_, new_n6187_, new_n10873_, new_n6188_, new_n10885_,
    new_n6189_, new_n7445_, new_n10893_, new_n6190_, new_n10906_,
    new_n6191_, new_n10914_, new_n6192_, new_n10927_, new_n6193_,
    new_n10935_, new_n6194_, new_n7446_, new_n10948_, new_n6195_,
    new_n10957_, new_n6196_, new_n10967_, new_n6197_, new_n10975_,
    new_n6198_, new_n10984_, new_n6199_, new_n7845_, new_n10992_,
    new_n6200_, new_n11000_, new_n6201_, new_n11008_, new_n6202_,
    new_n11047_, new_n6203_, new_n11075_, new_n6204_, new_n7027_,
    new_n7066_, new_n7447_, new_n11076_, new_n6205_, new_n6206_,
    new_n11096_, new_n6207_, new_n11102_, new_n6208_, new_n11126_,
    new_n6209_, new_n11149_, new_n7448_, new_n6210_, new_n11169_,
    new_n6211_, new_n6212_, new_n11190_, new_n6213_, new_n11201_,
    new_n6214_, new_n11227_, new_n6215_, new_n7449_, new_n11228_,
    new_n6216_, new_n11239_, new_n6217_, new_n11265_, new_n6218_,
    new_n11266_, new_n6219_, new_n11277_, new_n6220_, new_n7450_,
    new_n6221_, new_n11340_, new_n6222_, new_n11308_, new_n6223_,
    new_n11349_, new_n6224_, new_n11361_, new_n6225_, new_n11378_,
    new_n9540_, new_n6226_, new_n11384_, new_n6227_, new_n11388_,
    new_n6228_, new_n11404_, new_n6229_, new_n11414_, new_n6230_,
    new_n11424_, new_n7451_, new_n6231_, new_n11445_, new_n6232_,
    new_n11450_, new_n6233_, new_n11454_, new_n6234_, new_n11468_,
    new_n6235_, new_n7802_, new_n7452_, new_n6236_, new_n6237_, new_n7822_,
    new_n6238_, new_n6239_, new_n7839_, new_n6240_, new_n6241_, new_n7856_,
    new_n6242_, new_n7453_, new_n6243_, new_n7873_, new_n6244_, new_n6245_,
    new_n7890_, new_n6246_, new_n6247_, new_n7907_, new_n6248_, new_n6249_,
    new_n7879_, new_n7924_, new_n6250_, new_n6251_, new_n7941_, new_n6252_,
    new_n6253_, new_n7958_, new_n6254_, new_n6255_, new_n7975_, new_n7454_,
    new_n6256_, new_n6257_, new_n7992_, new_n6258_, new_n6259_, new_n8009_,
    new_n6260_, new_n6261_, new_n8026_, new_n6262_, new_n10478_,
    new_n7455_, new_n6263_, new_n8043_, new_n6264_, new_n6265_, new_n8060_,
    new_n6266_, new_n6267_, new_n8077_, new_n6268_, new_n6269_, new_n7456_,
    new_n8094_, new_n6270_, new_n6271_, new_n8111_, new_n6272_, new_n6273_,
    new_n8130_, new_n6274_, new_n6275_, new_n8147_, new_n7828_, new_n6276_,
    new_n6277_, new_n8165_, new_n6278_, new_n6279_, new_n8182_, new_n6280_,
    new_n6281_, new_n8200_, new_n6282_, new_n7457_, new_n6283_, new_n6284_,
    new_n8233_, new_n6285_, new_n6286_, new_n8250_, new_n6287_, new_n6288_,
    new_n8268_, new_n6289_, new_n7458_, new_n6290_, new_n8437_, new_n6291_,
    new_n10430_, new_n6292_, new_n10434_, new_n6293_, new_n6294_,
    new_n10439_, new_n6295_, new_n7459_, new_n10443_, new_n6296_,
    new_n10450_, new_n6297_, new_n10453_, new_n6298_, new_n6299_,
    new_n10458_, new_n6300_, new_n10462_, new_n7460_, new_n6301_,
    new_n6302_, new_n6303_, new_n10582_, new_n6304_, new_n10599_,
    new_n6305_, new_n10620_, new_n6306_, new_n10632_, new_n7461_,
    new_n6307_, new_n6308_, new_n10655_, new_n6309_, new_n10681_,
    new_n6310_, new_n7588_, new_n6311_, new_n7602_, new_n6312_, new_n8415_,
    new_n7627_, new_n6313_, new_n7641_, new_n6314_, new_n7670_, new_n6315_,
    new_n7685_, new_n6316_, new_n7740_, new_n6317_, new_n7462_, new_n8405_,
    new_n6318_, new_n6319_, new_n6320_, new_n8493_, new_n6321_, new_n6322_,
    new_n6323_, new_n6324_, new_n6325_, new_n7067_, new_n7463_, new_n8725_,
    new_n6326_, new_n8730_, new_n6327_, new_n6328_, new_n8798_, new_n6329_,
    new_n6330_, new_n8839_, new_n6331_, new_n7464_, new_n6332_, new_n6333_,
    new_n9099_, new_n6334_, new_n9164_, new_n6335_, new_n9562_, new_n6336_,
    new_n9566_, new_n6337_, new_n7465_, new_n9552_, new_n6338_, new_n9631_,
    new_n6339_, new_n9735_, new_n6340_, new_n9812_, new_n6341_, new_n9904_,
    new_n6342_, new_n7466_, new_n10031_, new_n6343_, new_n10107_,
    new_n6344_, new_n10108_, new_n6345_, new_n10115_, new_n6346_,
    new_n10183_, new_n6347_, new_n7467_, new_n10497_, new_n6348_,
    new_n10509_, new_n6349_, new_n10520_, new_n6350_, new_n6351_,
    new_n6352_, new_n10587_, new_n6353_, new_n7468_, new_n10699_,
    new_n6354_, new_n6355_, new_n6356_, new_n6357_, new_n6358_, new_n6359_,
    new_n6360_, new_n6361_, new_n6362_, new_n7469_, new_n11057_,
    new_n6363_, new_n11071_, new_n6364_, new_n11091_, new_n6365_,
    new_n11143_, new_n6366_, new_n11164_, new_n6367_, new_n7470_,
    new_n11185_, new_n6368_, new_n11211_, new_n6369_, new_n11223_,
    new_n6370_, new_n11249_, new_n6371_, new_n11261_, new_n6372_,
    new_n9061_, new_n11288_, new_n6373_, new_n11301_, new_n6374_,
    new_n11372_, new_n6375_, new_n11396_, new_n6376_, new_n11408_,
    new_n6377_, new_n7471_, new_n11435_, new_n6378_, new_n6379_,
    new_n6380_, new_n6381_, new_n6382_, new_n10519_, new_n6383_,
    new_n10605_, new_n6384_, new_n10384_, new_n7472_, new_n10634_,
    new_n6385_, new_n10637_, new_n6386_, new_n6387_, new_n6388_,
    new_n6389_, new_n6390_, new_n6391_, new_n6392_, new_n7473_, new_n6393_,
    new_n6394_, new_n6395_, new_n6396_, new_n6397_, new_n6398_, new_n6399_,
    new_n6400_, new_n6401_, new_n10881_, new_n7474_, new_n6402_,
    new_n6403_, new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_,
    new_n6409_, new_n6410_, new_n6411_, new_n9003_, new_n6412_, new_n6413_,
    new_n6414_, new_n6415_, new_n6416_, new_n6417_, new_n8672_, new_n6418_,
    new_n9191_, new_n6419_, new_n7475_, new_n9281_, new_n6420_, new_n9284_,
    new_n6421_, new_n6422_, new_n10606_, new_n6423_, new_n6424_,
    new_n6425_, new_n6426_, new_n10407_, new_n6427_, new_n6428_,
    new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_, new_n6434_,
    new_n6435_, new_n6436_, new_n7476_, new_n6437_, new_n6438_, new_n6439_,
    new_n10883_, new_n6440_, new_n6441_, new_n6442_, new_n6443_,
    new_n6444_, new_n6445_, new_n8533_, new_n6446_, new_n6447_, new_n6448_,
    new_n6449_, new_n6450_, new_n6451_, new_n6452_, new_n6453_, new_n6454_,
    new_n6455_, new_n7477_, new_n6456_, new_n7736_, new_n6457_, new_n7789_,
    new_n6458_, new_n7796_, new_n6459_, new_n8287_, new_n6460_, new_n6461_,
    new_n7478_, new_n8465_, new_n6462_, new_n8477_, new_n6463_, new_n8507_,
    new_n6464_, new_n6465_, new_n8530_, new_n6466_, new_n8540_, new_n7068_,
    new_n7479_, new_n6467_, new_n8545_, new_n6468_, new_n8547_, new_n6469_,
    new_n8562_, new_n6470_, new_n8568_, new_n6471_, new_n8581_, new_n7480_,
    new_n6472_, new_n8590_, new_n6473_, new_n8607_, new_n6474_, new_n8633_,
    new_n6475_, new_n8648_, new_n6476_, new_n8656_, new_n7481_, new_n6477_,
    new_n8663_, new_n6478_, new_n8683_, new_n6479_, new_n8689_, new_n6480_,
    new_n8692_, new_n6481_, new_n8707_, new_n7482_, new_n6482_, new_n8718_,
    new_n6483_, new_n8723_, new_n6484_, new_n8740_, new_n6485_, new_n8746_,
    new_n6486_, new_n8759_, new_n7483_, new_n6487_, new_n8766_, new_n6488_,
    new_n8786_, new_n6489_, new_n8793_, new_n6490_, new_n8796_, new_n6491_,
    new_n8814_, new_n7484_, new_n6492_, new_n6493_, new_n8829_, new_n6494_,
    new_n8837_, new_n6495_, new_n8851_, new_n6496_, new_n8861_, new_n6497_,
    new_n10377_, new_n8878_, new_n6498_, new_n8884_, new_n6499_,
    new_n8897_, new_n6500_, new_n8908_, new_n6501_, new_n8915_, new_n6502_,
    new_n7485_, new_n8918_, new_n6503_, new_n6504_, new_n8937_, new_n6505_,
    new_n8946_, new_n6506_, new_n8961_, new_n6507_, new_n6508_, new_n7486_,
    new_n8976_, new_n6509_, new_n8987_, new_n6510_, new_n6511_, new_n9010_,
    new_n6512_, new_n9015_, new_n6513_, new_n6514_, new_n7487_, new_n9034_,
    new_n6515_, new_n9040_, new_n6516_, new_n9052_, new_n6517_, new_n6518_,
    new_n9067_, new_n6519_, new_n9087_, new_n9280_, new_n7586_, new_n6520_,
    new_n9095_, new_n6521_, new_n9097_, new_n6522_, new_n9115_, new_n6523_,
    new_n6524_, new_n9130_, new_n6525_, new_n7488_, new_n6526_, new_n6527_,
    new_n9160_, new_n6528_, new_n9162_, new_n6529_, new_n9182_, new_n6530_,
    new_n9189_, new_n6531_, new_n7489_, new_n9205_, new_n6532_, new_n9212_,
    new_n6533_, new_n9225_, new_n6534_, new_n9232_, new_n6535_, new_n9238_,
    new_n6536_, new_n7490_, new_n9253_, new_n6537_, new_n9260_, new_n6538_,
    new_n6539_, new_n6540_, new_n9318_, new_n6541_, new_n6542_, new_n6543_,
    new_n7491_, new_n9342_, new_n6544_, new_n6545_, new_n6546_, new_n9365_,
    new_n6547_, new_n6548_, new_n9380_, new_n6549_, new_n6550_, new_n7492_,
    new_n6551_, new_n6552_, new_n6553_, new_n6554_, new_n9423_, new_n6555_,
    new_n6556_, new_n9438_, new_n6557_, new_n6558_, new_n7493_, new_n9453_,
    new_n6559_, new_n6560_, new_n9468_, new_n6561_, new_n6562_, new_n9482_,
    new_n6563_, new_n6564_, new_n9498_, new_n7494_, new_n6565_, new_n6566_,
    new_n6567_, new_n9520_, new_n6568_, new_n6569_, new_n9578_, new_n6570_,
    new_n9592_, new_n6571_, new_n7495_, new_n9607_, new_n6572_, new_n9622_,
    new_n6573_, new_n9636_, new_n6574_, new_n9639_, new_n6575_, new_n9657_,
    new_n6576_, new_n7496_, new_n9672_, new_n6577_, new_n9697_, new_n6578_,
    new_n9707_, new_n6579_, new_n9720_, new_n6580_, new_n9758_, new_n6581_,
    new_n7069_, new_n7497_, new_n9772_, new_n6582_, new_n9786_, new_n6583_,
    new_n9800_, new_n6584_, new_n9833_, new_n6585_, new_n9848_, new_n6586_,
    new_n7498_, new_n9863_, new_n6587_, new_n9885_, new_n6588_, new_n9896_,
    new_n6589_, new_n6590_, new_n9922_, new_n6591_, new_n6592_, new_n7499_,
    new_n9942_, new_n6593_, new_n9956_, new_n6594_, new_n9967_, new_n6595_,
    new_n9982_, new_n6596_, new_n9996_, new_n6597_, new_n7500_, new_n9999_,
    new_n6598_, new_n10001_, new_n6599_, new_n10040_, new_n6600_,
    new_n10048_, new_n6601_, new_n6602_, new_n10061_, new_n7501_,
    new_n6603_, new_n10125_, new_n6604_, new_n6605_, new_n10169_,
    new_n6606_, new_n10176_, new_n6607_, new_n10182_, new_n6608_,
    new_n7502_, new_n10192_, new_n6609_, new_n10321_, new_n6610_,
    new_n10331_, new_n6611_, new_n6612_, new_n6613_, new_n10514_,
    new_n6614_, new_n7503_, new_n10518_, new_n6615_, new_n6616_,
    new_n10636_, new_n6617_, new_n10666_, new_n6618_, new_n10688_,
    new_n6619_, new_n10696_, new_n7504_, new_n6620_, new_n10711_,
    new_n6621_, new_n10720_, new_n6622_, new_n11031_, new_n6623_,
    new_n11108_, new_n6624_, new_n11113_, new_n7505_, new_n6625_,
    new_n11119_, new_n6626_, new_n11123_, new_n6627_, new_n11148_,
    new_n6628_, new_n11306_, new_n6629_, new_n11360_, new_n7506_,
    new_n6630_, new_n11363_, new_n6631_, new_n11377_, new_n6632_,
    new_n11399_, new_n6633_, new_n11403_, new_n6634_, new_n11437_,
    new_n8515_, new_n7507_, new_n6635_, new_n11444_, new_n6636_,
    new_n11449_, new_n6637_, new_n11453_, new_n6638_, new_n11463_,
    new_n6639_, new_n11467_, new_n7508_, new_n6640_, new_n6641_,
    new_n6642_, new_n6643_, new_n6644_, new_n6645_, new_n6646_, new_n6647_,
    new_n6648_, new_n6649_, new_n7930_, new_n6650_, new_n6651_, new_n6652_,
    new_n6653_, new_n6654_, new_n6655_, new_n6656_, new_n6657_, new_n6658_,
    new_n6659_, new_n7509_, new_n6660_, new_n6661_, new_n6662_, new_n6663_,
    new_n6664_, new_n6665_, new_n6666_, new_n6667_, new_n6668_, new_n6669_,
    new_n7510_, new_n6670_, new_n6671_, new_n6672_, new_n6673_, new_n6674_,
    new_n6675_, new_n6676_, new_n6677_, new_n6678_, new_n6679_, new_n7511_,
    new_n6680_, new_n6681_, new_n6682_, new_n6683_, new_n6684_, new_n6685_,
    new_n6686_, new_n6687_, new_n6688_, new_n6689_, new_n7862_, new_n6690_,
    new_n6691_, new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_,
    new_n8412_, new_n6697_, new_n6698_, new_n7512_, new_n8438_, new_n6699_,
    new_n6700_, new_n6701_, new_n6702_, new_n6703_, new_n10431_,
    new_n6704_, new_n10435_, new_n6705_, new_n7513_, new_n10444_,
    new_n6706_, new_n6707_, new_n10451_, new_n6708_, new_n10459_,
    new_n6709_, new_n6710_, new_n10486_, new_n6711_, new_n7514_,
    new_n6712_, new_n10537_, new_n6713_, new_n6714_, new_n10600_,
    new_n6715_, new_n6716_, new_n6717_, new_n6718_, new_n10682_,
    new_n7070_, new_n7515_, new_n6719_, new_n6720_, new_n6721_, new_n6722_,
    new_n6723_, new_n6724_, new_n6725_, new_n6726_, new_n6727_, new_n6728_,
    new_n7516_, new_n6729_, new_n6730_, new_n6731_, new_n6732_, new_n6733_,
    new_n6734_, new_n6735_, new_n8288_, new_n6736_, new_n6737_, new_n7517_,
    new_n6738_, new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_,
    new_n6744_, new_n6745_, new_n6746_, new_n6747_, new_n7518_, new_n6748_,
    new_n6749_, new_n6750_, new_n6751_, new_n6752_, new_n6753_, new_n6754_,
    new_n6755_, new_n6756_, new_n6757_, new_n7519_, new_n6758_, new_n6759_,
    new_n6760_, new_n6761_, new_n6762_, new_n6763_, new_n6764_, new_n6765_,
    new_n6766_, new_n6767_, new_n7808_, new_n6768_, new_n6769_, new_n6770_,
    new_n6771_, new_n6772_, new_n6773_, new_n6774_, new_n9279_, new_n6775_,
    new_n9304_, new_n9125_, new_n6776_, new_n9539_, new_n6777_, new_n9542_,
    new_n6778_, new_n6779_, new_n6780_, new_n9585_, new_n6781_, new_n6782_,
    new_n7520_, new_n9614_, new_n6783_, new_n6784_, new_n6785_, new_n9650_,
    new_n6786_, new_n6787_, new_n9699_, new_n6788_, new_n6789_, new_n7521_,
    new_n6790_, new_n6791_, new_n6792_, new_n9750_, new_n6793_, new_n6794_,
    new_n9779_, new_n6795_, new_n9792_, new_n6796_, new_n7522_, new_n9806_,
    new_n6797_, new_n6798_, new_n6799_, new_n6800_, new_n9840_, new_n6801_,
    new_n9855_, new_n6802_, new_n6803_, new_n7071_, new_n10412_,
    new_n6804_, new_n9889_, new_n6805_, new_n6806_, new_n6807_, new_n9929_,
    new_n6808_, new_n6809_, new_n9960_, new_n6810_, new_n7523_, new_n9974_,
    new_n6811_, new_n6812_, new_n6813_, new_n10103_, new_n6814_,
    new_n6815_, new_n6816_, new_n6817_, new_n10403_, new_n7524_,
    new_n6818_, new_n6819_, new_n10507_, new_n6820_, new_n10541_,
    new_n6821_, new_n10562_, new_n6822_, new_n6823_, new_n6824_,
    new_n7525_, new_n10701_, new_n6825_, new_n6826_, new_n6827_,
    new_n6828_, new_n11020_, new_n6829_, new_n11023_, new_n6830_,
    new_n6831_, new_n7526_, new_n6832_, new_n6833_, new_n11082_,
    new_n6834_, new_n6835_, new_n6836_, new_n6837_, new_n6838_, new_n6839_,
    new_n6840_, new_n7527_, new_n6841_, new_n6842_, new_n6843_, new_n6844_,
    new_n6845_, new_n6846_, new_n6847_, new_n6848_, new_n6849_, new_n6850_,
    new_n7528_, new_n6851_, new_n6852_, new_n6853_, new_n6854_, new_n6855_,
    new_n6856_, new_n6857_, new_n6858_, new_n6859_, new_n6860_, new_n7529_,
    new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_, new_n6866_,
    new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n7530_, new_n6871_,
    new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_,
    new_n6878_, new_n6879_, new_n6880_, new_n7531_, new_n6881_, new_n6882_,
    new_n6883_, new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_,
    new_n6889_, new_n6890_, new_n7028_, new_n7072_, new_n7532_, new_n6891_,
    new_n6892_, new_n6893_, new_n6894_, new_n6895_, new_n6896_, new_n6897_,
    new_n6898_, new_n6899_, new_n6900_, new_n7533_, new_n6901_, new_n6902_,
    new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_, new_n6908_,
    new_n6909_, new_n6910_, new_n7534_, new_n9906_, new_n6911_, new_n6912_,
    new_n6913_, new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_,
    new_n10117_, new_n7535_, new_n6919_, new_n10282_, new_n6920_,
    new_n6921_, new_n10398_, new_n6922_, new_n6923_, new_n10506_,
    new_n6924_, new_n6925_, new_n7536_, new_n10568_, new_n6926_,
    new_n6927_, new_n10561_, new_n6928_, new_n6929_, new_n6930_,
    new_n11010_, new_n6931_, new_n11024_, new_n7537_, new_n6932_,
    new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_, new_n6938_,
    new_n6939_, new_n6940_, new_n6941_, new_n7538_, new_n6942_, new_n6943_,
    new_n6944_, new_n6945_, new_n8888_, new_n6946_, new_n6947_, new_n9709_,
    new_n6948_, new_n9722_, new_n7896_, new_n6949_, new_n9774_, new_n6950_,
    new_n9958_, new_n6951_, new_n6952_, new_n10739_, new_n6953_,
    new_n10965_, new_n6954_, new_n7539_, new_n6955_, new_n8939_,
    new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_,
    new_n6962_, new_n6963_, new_n7540_, new_n6964_, new_n6965_, new_n6966_,
    new_n6967_, new_n6968_, new_n6969_, new_n6970_, new_n9624_, new_n6971_,
    new_n9760_, new_n7073_, new_n7541_, new_n6972_, new_n9788_, new_n6973_,
    new_n9802_, new_n6974_, new_n9887_, new_n6975_, new_n9984_, new_n6976_,
    new_n6977_, new_n7542_, new_n6978_, new_n6979_, new_n6980_, new_n6981_,
    new_n6982_, new_n6983_, new_n6984_, new_n6985_, new_n6986_, new_n6987_,
    new_n7543_, new_n6988_, new_n6989_, new_n6990_, new_n6991_, new_n6992_,
    new_n6993_, new_n6994_, new_n11103_, new_n6995_, new_n10324_,
    new_n7544_, new_n6996_, new_n6997_, new_n6998_, new_n11294_,
    new_n6999_, new_n11447_, new_n7000_, new_n11432_, new_n7001_,
    new_n11428_, new_n7545_, new_n7002_, new_n7003_, new_n7004_,
    new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_, new_n7010_,
    new_n7011_, new_n7546_, new_n7012_, new_n7013_, new_n7014_, new_n7015_,
    new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_,
    new_n7547_, new_n8865_, new_n7548_, new_n7549_, new_n7550_, new_n7074_,
    new_n7551_, new_n7552_, new_n9313_, new_n7553_, new_n9311_, new_n7554_,
    new_n7555_, new_n7556_, new_n7557_, new_n7558_, new_n7075_, new_n7559_,
    new_n7809_, new_n7560_, new_n7561_, new_n7562_, new_n7563_, new_n7564_,
    new_n7565_, new_n7566_, new_n9299_, new_n7567_, new_n7568_, new_n7569_,
    new_n7579_, new_n7585_, new_n7582_, new_n7584_, new_n7600_, new_n7076_,
    new_n7599_, new_n7607_, new_n7601_, new_n7620_, new_n7625_, new_n7622_,
    new_n7624_, new_n7639_, new_n7077_, new_n7637_, new_n7642_, new_n7649_,
    new_n7650_, new_n7661_, new_n7663_, new_n7668_, new_n7666_, new_n7671_,
    new_n11230_, new_n7682_, new_n7680_, new_n7686_, new_n7693_,
    new_n7694_, new_n7705_, new_n7707_, new_n7712_, new_n7078_, new_n7684_,
    new_n7715_, new_n7669_, new_n7718_, new_n7640_, new_n7732_, new_n7729_,
    new_n7735_, new_n7737_, new_n7734_, new_n7079_, new_n7710_, new_n7741_,
    new_n7688_, new_n7744_, new_n7672_, new_n7747_, new_n7644_, new_n7750_,
    new_n7754_, new_n7753_, new_n7029_, new_n11078_, new_n7758_,
    new_n7757_, new_n7762_, new_n7761_, new_n7765_, new_n7781_, new_n7786_,
    new_n7080_, new_n7788_, new_n8406_, new_n7081_, new_n8114_, new_n8150_,
    new_n8185_, new_n8220_, new_n8449_, new_n8217_, new_n8253_, new_n8284_,
    new_n8286_, new_n8289_, new_n7814_, new_n7082_, new_n8508_, new_n7083_,
    new_n8569_, new_n8402_, new_n7775_, new_n8414_, new_n8310_, new_n7799_,
    new_n7084_, new_n7794_, new_n8455_, new_n8313_, new_n8466_, new_n8470_,
    new_n7806_, new_n8479_, new_n7807_, new_n8481_, new_n7030_, new_n8634_,
    new_n8316_, new_n8491_, new_n8494_, new_n8498_, new_n8501_, new_n7826_,
    new_n7827_, new_n8511_, new_n8516_, new_n7085_, new_n8319_, new_n8531_,
    new_n7843_, new_n8542_, new_n7844_, new_n8546_, new_n8544_, new_n8322_,
    new_n7086_, new_n8563_, new_n7860_, new_n7861_, new_n8325_, new_n8582_,
    new_n8583_, new_n7877_, new_n8592_, new_n7878_, new_n7087_, new_n8597_,
    new_n8328_, new_n8608_, new_n8611_, new_n8625_, new_n7894_, new_n7895_,
    new_n8635_, new_n7088_, new_n8331_, new_n8649_, new_n7911_, new_n8658_,
    new_n7912_, new_n8664_, new_n8668_, new_n8665_, new_n8334_, new_n7089_,
    new_n8684_, new_n8652_, new_n7928_, new_n8693_, new_n8694_, new_n8337_,
    new_n8708_, new_n7945_, new_n8724_, new_n7090_, new_n8673_, new_n8727_,
    new_n8340_, new_n8741_, new_n7962_, new_n7963_, new_n8343_, new_n8760_,
    new_n8503_, new_n7979_, new_n7980_, new_n8775_, new_n8770_, new_n8346_,
    new_n8787_, new_n7996_, new_n7997_, new_n8797_, new_n7091_, new_n8795_,
    new_n8349_, new_n8013_, new_n8014_, new_n8834_, new_n8838_, new_n8352_,
    new_n8852_, new_n10810_, new_n8030_, new_n8031_, new_n8355_,
    new_n8879_, new_n8047_, new_n8048_, new_n8889_, new_n8894_, new_n8898_;
  
  
// BEGIN WF
parameter WF_N = 16;     // TOKEN_N // set by python
parameter WF_DEPTH = 6; // TOKEN_STAGES // set by python
parameter LOCKABLE_INPUTS = 16;  // TOKEN_WF_LOCKABLE_INPUTS modify 32 to be whatever your total lockable bits are
// END WF

// WF BEGIN
// TOKEN_CORRECT_KEYS
// correct key0: 48'b110101010010111001110101001010010010000101001101
// correct key1: 48'b011111101011111000001000011101011111000010100000
// correct key2: 48'b001010010001101010111111001100010111011000111111
input [3*WF_N*WF_DEPTH/2-1:0] keyinput;
wire   [WF_N*WF_DEPTH/2-1:0]  key0;
wire   [WF_N*WF_DEPTH/2-1:0]  key1;
wire   [WF_N*WF_DEPTH/2-1:0]  key2;

wire [LOCKABLE_INPUTS-1:0] addressable_wf_inputs;
wire [WF_N-1:0] wf_inputs;
wire [WF_N-1:0] wf_outputs;
wire [LOCKABLE_INPUTS-1:0] addressable_wf_outputs;

// modify these to be the locked versions of the wires you're locking

//wire [7:0] input1_wflocked;         // 8 wide
//wire [7:0] input2_wflocked;         // 8 wide
// WF END

wire new_n10564_in, new_n8671_in, new_n11341_in, new_n10479_in,
      new_n10426_in, new_n10006_in, new_n10209_in, new_n10034_in,
      new_n10196_in, new_n9544_in, new_n8670_in, new_n8519_in,
      new_n7725_in, new_n10487_in, new_n10621_in, new_n7137_in;

// WF BEGIN

assign key0 = keyinput[WF_N*WF_DEPTH/2-1:0];
assign key1 = keyinput[WF_N*WF_DEPTH-1:WF_N*WF_DEPTH/2];
assign key2 = keyinput[3*WF_N*WF_DEPTH/2-1:WF_N*WF_DEPTH];

assign addressable_wf_inputs = {  // length must match LOCKABLE_INPUTS
  new_n10564_in, new_n8671_in, new_n11341_in, new_n10479_in,
  new_n10426_in, new_n10006_in, new_n10209_in, new_n10034_in,
  new_n10196_in, new_n9544_in, new_n8670_in, new_n8519_in,
  new_n7725_in, new_n10487_in, new_n10621_in, new_n7137_in  // modify this to whatever wires you want to lock
};

//for up to N = LOCKABLE_INPUTS rounded down to nearest even number
// TOKEN_PICK_WF_INPUTS
//assign addressable_wf_outputs[15] = addressable_wf_inputs[15];
//assign addressable_wf_outputs[14] = addressable_wf_inputs[14];
//assign addressable_wf_outputs[13] = addressable_wf_inputs[13];
//assign addressable_wf_outputs[12] = addressable_wf_inputs[12];
//assign addressable_wf_outputs[11] = addressable_wf_inputs[11];
//assign addressable_wf_outputs[10] = addressable_wf_inputs[10];
//assign addressable_wf_outputs[9] = addressable_wf_inputs[9];
//assign addressable_wf_outputs[8] = addressable_wf_inputs[8];
//assign addressable_wf_outputs[7] = addressable_wf_inputs[7];
//assign addressable_wf_outputs[6] = addressable_wf_inputs[6];
//assign addressable_wf_outputs[5] = addressable_wf_inputs[5];
//assign addressable_wf_outputs[4] = addressable_wf_inputs[4];
//assign addressable_wf_outputs[3] = addressable_wf_inputs[3];
//assign addressable_wf_outputs[2] = addressable_wf_inputs[2];
//assign addressable_wf_outputs[1] = addressable_wf_inputs[1];
//assign addressable_wf_outputs[0] = addressable_wf_inputs[0];


// TOKEN_BEGIN_WF_IN_ASSIGN
assign wf_inputs[15] = addressable_wf_inputs[12];
assign wf_inputs[14] = addressable_wf_inputs[0];
assign wf_inputs[13] = addressable_wf_inputs[10];
assign wf_inputs[12] = addressable_wf_inputs[8];
assign wf_inputs[11] = addressable_wf_inputs[9];
assign wf_inputs[10] = addressable_wf_inputs[13];
assign wf_inputs[9] = addressable_wf_inputs[5];
assign wf_inputs[8] = addressable_wf_inputs[3];
assign wf_inputs[7] = addressable_wf_inputs[11];
assign wf_inputs[6] = addressable_wf_inputs[7];
assign wf_inputs[5] = addressable_wf_inputs[2];
assign wf_inputs[4] = addressable_wf_inputs[4];
assign wf_inputs[3] = addressable_wf_inputs[1];
assign wf_inputs[2] = addressable_wf_inputs[14];
assign wf_inputs[1] = addressable_wf_inputs[15];
assign wf_inputs[0] = addressable_wf_inputs[6];


wf_8x6 #(.N(WF_N), .stages(WF_DEPTH)) wf0 (  // TOKEN_WF_MODNAME
.IN(wf_inputs),
.K0(key0),
.K1(key1),
.K2(key2),
.OUT(wf_outputs)
);

// TOKEN_BEGIN_WF_OUT_ASSIGN
assign addressable_wf_outputs[12] = wf_outputs[15];
assign addressable_wf_outputs[0] = wf_outputs[14];
assign addressable_wf_outputs[10] = wf_outputs[13];
assign addressable_wf_outputs[8] = wf_outputs[12];
assign addressable_wf_outputs[9] = wf_outputs[11];
assign addressable_wf_outputs[13] = wf_outputs[10];
assign addressable_wf_outputs[5] = wf_outputs[9];
assign addressable_wf_outputs[3] = wf_outputs[8];
assign addressable_wf_outputs[11] = wf_outputs[7];
assign addressable_wf_outputs[7] = wf_outputs[6];
assign addressable_wf_outputs[2] = wf_outputs[5];
assign addressable_wf_outputs[4] = wf_outputs[4];
assign addressable_wf_outputs[1] = wf_outputs[3];
assign addressable_wf_outputs[14] = wf_outputs[2];
assign addressable_wf_outputs[15] = wf_outputs[1];
assign addressable_wf_outputs[6] = wf_outputs[0];


assign new_n10564_ = addressable_wf_outputs[15];
assign new_n8671_ = addressable_wf_outputs[14];
assign new_n11341_ = addressable_wf_outputs[13];
assign new_n10479_ = addressable_wf_outputs[12];
assign new_n10426_ = addressable_wf_outputs[11];
assign new_n10006_ = addressable_wf_outputs[10];
assign new_n10209_ = addressable_wf_outputs[9];
assign new_n10034_ = addressable_wf_outputs[8];
assign new_n10196_ = addressable_wf_outputs[7];
assign new_n9544_ = addressable_wf_outputs[6];
assign new_n8670_ = addressable_wf_outputs[5];
assign new_n8519_ = addressable_wf_outputs[4];
assign new_n7725_ = addressable_wf_outputs[3];
assign new_n10487_ = addressable_wf_outputs[2];
assign new_n10621_ = addressable_wf_outputs[1];
assign new_n7137_ = addressable_wf_outputs[0];
//assign input1_wflocked = addressable_wf_outputs[7:0];  // modify these to be whatever wires are locked
//assign input2_wflocked = addressable_wf_outputs[15:8];  // modify these to be whatever wires are locked
// Don't forget to replace original wires with wflocked variants
// WF END
  
  
  assign new_n7022_ = ~new_n8865_;
  assign new_n7031_ = ~new_n8214_;
  assign new_n7092_ = ~new_n10810_;
  assign n559 = ~new_n6101_ | ~new_n5807_;
  assign new_n8358_ = new_n6875_ | new_n6757_;
  assign new_n8909_ = new_n8910_ ^ new_n8911_;
  assign new_n8064_ = ~new_n8916_ ^ new_n8066_;
  assign new_n8065_ = new_n8917_ & new_n6503_;
  assign new_n8919_ = new_n8920_ & new_n6504_;
  assign new_n8920_ = new_n7436_ | new_n7518_;
  assign new_n8917_ = new_n7113_ | new_n6758_;
  assign n554 = ~new_n6102_ | ~new_n5808_;
  assign new_n8361_ = new_n6876_ | new_n6759_;
  assign new_n7093_ = ~new_n7629_;
  assign new_n8938_ = new_n6956_ ^ new_n8940_;
  assign new_n8081_ = new_n6333_ & new_n7090_;
  assign new_n8082_ = new_n7436_ ^ new_n8940_;
  assign n549 = ~new_n6105_ | ~new_n5810_;
  assign new_n8364_ = new_n6877_ | new_n6760_;
  assign new_n8098_ = ~new_n8117_ ^ new_n8100_;
  assign new_n8099_ = ~new_n7336_ ^ new_n8971_;
  assign new_n8979_ = new_n7117_ & new_n7337_;
  assign new_n8984_ = new_n7182_ & new_n6510_;
  assign new_n8988_ = new_n9043_ & new_n8989_;
  assign new_n8548_ = new_n7240_ & new_n7512_;
  assign n544 = ~new_n6107_ | ~new_n5812_;
  assign new_n8367_ = new_n6878_ | new_n6761_;
  assign new_n9001_ = new_n7211_ | new_n8968_;
  assign new_n9011_ = new_n7181_ & new_n7266_;
  assign new_n8118_ = new_n9014_ & new_n6513_;
  assign new_n9016_ = new_n9017_ & new_n6514_;
  assign new_n9017_ = new_n7433_ | new_n7535_;
  assign new_n9014_ = new_n7114_ | new_n6762_;
  assign n539 = ~new_n6108_ | ~new_n5813_;
  assign new_n8370_ = new_n6879_ | new_n6763_;
  assign new_n7094_ = ~new_n8548_;
  assign new_n9035_ = ~new_n7428_ ^ new_n7366_;
  assign new_n8134_ = ~new_n8152_ ^ new_n8136_;
  assign new_n8135_ = ~new_n7433_ ^ new_n7428_;
  assign n534 = ~new_n6111_ | ~new_n5815_;
  assign new_n8373_ = new_n6880_ | new_n6764_;
  assign new_n9063_ = new_n9059_ | new_n7372_;
  assign new_n9068_ = new_n7183_ & new_n7267_;
  assign new_n8153_ = ~new_n7337_ ^ new_n9057_;
  assign new_n9076_ = new_n7420_ | new_n7534_;
  assign new_n9071_ = new_n7218_ | new_n9101_;
  assign new_n7095_ = ~new_n9285_;
  assign n529 = ~new_n6112_ | ~new_n5818_;
  assign new_n8376_ = new_n6881_ | new_n6765_;
  assign new_n9088_ = ~new_n9089_ ^ new_n7372_;
  assign new_n8169_ = ~new_n8187_ ^ new_n8171_;
  assign new_n8170_ = new_n9096_ & new_n6522_;
  assign new_n9098_ = new_n6334_ & new_n7420_;
  assign new_n9096_ = new_n7218_ | new_n6766_;
  assign n524 = ~new_n6114_ | ~new_n5819_;
  assign new_n8379_ = new_n6882_ | new_n6767_;
  assign new_n9131_ = new_n7184_ & new_n7268_;
  assign new_n7096_ = ~new_n7628_;
  assign new_n8188_ = ~new_n7334_ ^ new_n9120_;
  assign new_n9136_ = new_n7219_ | new_n9166_;
  assign new_n9135_ = new_n9138_ & new_n6526_;
  assign new_n9138_ = new_n7421_ | new_n7533_;
  assign n519 = ~new_n6116_ | ~new_n5821_;
  assign new_n8382_ = new_n6883_ | new_n6768_;
  assign new_n9153_ = new_n7212_ | new_n9122_;
  assign new_n8204_ = ~new_n7429_ ^ new_n8206_;
  assign new_n8205_ = new_n9161_ & new_n6529_;
  assign new_n9163_ = new_n6335_ & new_n7421_;
  assign new_n9100_ = new_n7236_ & new_n7379_;
  assign new_n9161_ = new_n7219_ | new_n6769_;
  assign n514 = ~new_n6117_ | ~new_n5822_;
  assign new_n8385_ = new_n6884_ | new_n6770_;
  assign new_n9183_ = ~new_n9184_ ^ new_n7425_;
  assign new_n9190_ = new_n7185_ & new_n9133_;
  assign new_n9192_ = new_n7507_ | new_n8239_;
  assign new_n8223_ = ~new_n9166_ ^ new_n7425_;
  assign new_n9195_ = new_n7363_ | new_n8239_;
  assign n509 = ~new_n6118_ | ~new_n5823_;
  assign new_n8388_ = new_n6885_ | new_n6771_;
  assign new_n7097_ = ~new_n9100_;
  assign new_n9206_ = ~new_n9207_ ^ new_n9208_;
  assign new_n8237_ = ~new_n7507_ ^ new_n7531_;
  assign new_n8238_ = ~new_n7363_ ^ new_n9208_;
  assign n504 = ~new_n6119_ | ~new_n5825_;
  assign new_n8391_ = new_n6886_ | new_n6772_;
  assign new_n9226_ = ~new_n9227_ ^ new_n9228_;
  assign new_n9233_ = new_n7186_ & new_n7507_;
  assign new_n9234_ = new_n7394_ & new_n7549_;
  assign new_n9239_ = new_n7288_ & new_n7168_;
  assign n499 = ~new_n6120_ | ~new_n5826_;
  assign new_n10578_ = new_n10633_ & new_n7303_;
  assign new_n8394_ = new_n6887_ | new_n6773_;
  assign new_n8433_ = new_n9290_ & new_n9265_;
  assign new_n9254_ = new_n7506_ ^ new_n7427_;
  assign new_n8272_ = ~new_n7549_ ^ new_n9235_;
  assign new_n8273_ = ~new_n7427_ ^ new_n9243_;
  assign new_n9243_ = new_n9235_ & new_n10586_;
  assign n494 = ~new_n6123_ | ~new_n5827_;
  assign new_n8295_ = new_n9290_ & new_n7444_;
  assign new_n8292_ = new_n6888_ | new_n6774_;
  assign new_n9276_ = new_n7547_ | new_n6775_;
  assign new_n7098_ = ~new_n10578_;
  assign n489 = D_REG_31_ & new_n7567_;
  assign n484 = D_REG_30_ & new_n7567_;
  assign n479 = D_REG_29_ & new_n7567_;
  assign n474 = D_REG_28_ & new_n7567_;
  assign n469 = D_REG_27_ & new_n7567_;
  assign n464 = D_REG_26_ & new_n7567_;
  assign n459 = D_REG_25_ & new_n7567_;
  assign n454 = D_REG_24_ & new_n7567_;
  assign n449 = D_REG_23_ & new_n7567_;
  assign n444 = D_REG_22_ & new_n7567_;
  assign new_n7032_ = ~new_n8230_;
  assign new_n10172_ = new_n7290_ & new_n7280_;
  assign n439 = D_REG_21_ & new_n7567_;
  assign n434 = D_REG_20_ & new_n7567_;
  assign n429 = D_REG_19_ & new_n7567_;
  assign n424 = D_REG_18_ & new_n7567_;
  assign n419 = D_REG_17_ & new_n7567_;
  assign n414 = D_REG_16_ & new_n7567_;
  assign n409 = D_REG_15_ & new_n7567_;
  assign n404 = D_REG_14_ & new_n7567_;
  assign n399 = D_REG_13_ & new_n7567_;
  assign n394 = D_REG_12_ & new_n7567_;
  assign new_n7099_ = ~new_n10172_;
  assign n389 = D_REG_11_ & new_n7567_;
  assign n384 = D_REG_10_ & new_n7567_;
  assign n379 = D_REG_9_ & new_n7567_;
  assign n374 = D_REG_8_ & new_n7567_;
  assign n369 = D_REG_7_ & new_n7567_;
  assign n364 = D_REG_6_ & new_n7567_;
  assign n359 = D_REG_5_ & new_n7567_;
  assign n354 = D_REG_4_ & new_n7567_;
  assign n349 = D_REG_3_ & new_n7567_;
  assign n344 = D_REG_2_ & new_n7567_;
  assign new_n7100_ = ~new_n11017_;
  assign n339 = ~new_n6125_ | ~new_n5830_;
  assign n334 = ~new_n6126_ | ~new_n5831_;
  assign n329 = ~new_n6127_ | ~new_n9302_;
  assign new_n9302_ = new_n9303_ | new_n6776_;
  assign n324 = ~new_n9306_ | ~new_n5832_;
  assign new_n9312_ = new_n9303_ | new_n7552_;
  assign new_n9305_ = ~IR_REG_30_;
  assign new_n9314_ = new_n9313_ & new_n9303_;
  assign n319 = ~new_n9315_ | ~new_n5833_;
  assign new_n9319_ = new_n7162_ & new_n9303_;
  assign new_n8799_ = new_n7235_ & new_n7381_;
  assign new_n9303_ = new_n7297_ | IR_REG_29_;
  assign n314 = ~new_n9322_ | ~new_n5834_;
  assign n309 = ~new_n9330_ | ~new_n5836_;
  assign n304 = ~new_n9339_ | ~new_n5838_;
  assign n299 = ~new_n9344_ | ~new_n5839_;
  assign new_n9350_ = new_n7401_ & new_n9313_;
  assign n294 = ~new_n9353_ | ~new_n5841_;
  assign n289 = ~new_n9362_ | ~new_n5843_;
  assign new_n9366_ = new_n7165_ & new_n9359_;
  assign n284 = ~new_n9368_ | ~new_n5844_;
  assign new_n7101_ = ~new_n8799_;
  assign n279 = ~new_n9377_ | ~new_n5846_;
  assign new_n9381_ = new_n7164_ & new_n9374_;
  assign n274 = ~new_n9383_ | ~new_n5847_;
  assign n269 = ~new_n9392_ | ~new_n5849_;
  assign n264 = ~new_n9397_ | ~new_n5850_;
  assign n259 = ~new_n9406_ | ~new_n5852_;
  assign n254 = ~new_n9411_ | ~new_n5853_;
  assign n249 = ~new_n9420_ | ~new_n5855_;
  assign new_n9424_ = new_n9417_ & new_n7170_;
  assign n244 = ~new_n9426_ | ~new_n5856_;
  assign new_n9165_ = new_n7238_ & new_n7369_;
  assign n239 = ~new_n9435_ | ~new_n5858_;
  assign new_n9439_ = new_n9432_ & new_n7171_;
  assign n234 = ~new_n9441_ | ~new_n5859_;
  assign n229 = ~new_n9450_ | ~new_n5861_;
  assign new_n9454_ = new_n9447_ & new_n7172_;
  assign n224 = ~new_n9456_ | ~new_n5862_;
  assign n219 = ~new_n9465_ | ~new_n5864_;
  assign new_n9469_ = new_n7163_ & new_n9462_;
  assign n214 = ~new_n9471_ | ~new_n5865_;
  assign n209 = ~new_n9479_ | ~new_n5867_;
  assign new_n7102_ = ~new_n9165_;
  assign new_n9483_ = new_n7272_ & new_n7174_;
  assign n204 = ~new_n9486_ | ~new_n5868_;
  assign n199 = ~new_n9495_ | ~new_n5870_;
  assign n194 = ~new_n9500_ | ~new_n5871_;
  assign n189 = ~new_n9509_ | ~new_n5873_;
  assign n184 = ~new_n9517_ | ~new_n5875_;
  assign new_n9521_ = new_n7404_ & new_n7173_;
  assign n179 = ~new_n9524_ | ~new_n5876_;
  assign n174 = ~new_n6143_ | ~new_n5878_;
  assign n1337 = ~new_n9537_ | ~new_n9538_;
  assign new_n10521_ = new_n8257_ & new_n7257_;
  assign new_n9538_ = new_n10635_ | new_n6777_;
  assign n1327 = new_n6889_ | new_n6778_;
  assign new_n9549_ = new_n6338_ & new_n9553_;
  assign new_n9553_ = new_n7423_ | new_n6779_;
  assign new_n9558_ = new_n6336_ & new_n7412_;
  assign new_n9565_ = new_n6337_ & new_n7305_;
  assign n1322 = new_n6890_ | new_n6780_;
  assign new_n9579_ = ~new_n9580_ ^ new_n9581_;
  assign new_n9580_ = new_n7368_ ^ new_n9583_;
  assign n1317 = new_n6891_ | new_n6781_;
  assign new_n7103_ = ~new_n10521_;
  assign new_n9593_ = new_n9594_ ^ new_n9595_;
  assign new_n9594_ = ~new_n7222_ ^ new_n7376_;
  assign n1312 = new_n6892_ | new_n6782_;
  assign new_n9608_ = ~new_n9609_ ^ new_n9610_;
  assign new_n9610_ = ~new_n7360_ ^ new_n7374_;
  assign n1307 = new_n6893_ | new_n6783_;
  assign new_n9623_ = ~new_n9948_ ^ new_n6971_;
  assign n1302 = new_n6894_ | new_n6784_;
  assign new_n9629_ = new_n6339_ & new_n7199_;
  assign new_n9637_ = new_n9638_ & new_n6575_;
  assign new_n7774_ = new_n8406_ & new_n7772_;
  assign new_n9638_ = new_n7201_ | new_n6785_;
  assign n1297 = new_n6895_ | new_n6786_;
  assign new_n9658_ = new_n9659_ ^ new_n9660_;
  assign new_n9659_ = ~new_n9661_ ^ new_n9662_;
  assign n1292 = new_n6896_ | new_n6787_;
  assign new_n9673_ = new_n9674_ ^ new_n9675_;
  assign new_n9675_ = new_n6957_ ^ new_n6977_;
  assign new_n9674_ = ~new_n6947_ ^ new_n7569_;
  assign new_n9688_ = new_n7368_ | new_n9583_;
  assign new_n9581_ = new_n6958_ ^ new_n9685_;
  assign new_n7033_ = ~new_n9166_;
  assign new_n7104_ = ~new_n7774_;
  assign n1287 = new_n6897_ | new_n6788_;
  assign new_n9708_ = ~new_n6948_ ^ new_n7227_;
  assign n1282 = new_n6898_ | new_n6789_;
  assign new_n9721_ = ~new_n6949_ ^ new_n7228_;
  assign n1277 = new_n6899_ | new_n6790_;
  assign new_n9733_ = new_n6340_ & new_n9736_;
  assign new_n9736_ = new_n7423_ | new_n6791_;
  assign new_n9738_ = new_n7202_ | new_n6792_;
  assign n1272 = new_n6900_ | new_n6793_;
  assign new_n9759_ = ~new_n9905_ ^ new_n6972_;
  assign new_n7105_ = ~new_n8303_;
  assign n1267 = new_n6901_ | new_n6794_;
  assign new_n9773_ = ~new_n6950_ ^ new_n7345_;
  assign n1262 = new_n6902_ | new_n6795_;
  assign new_n9787_ = ~new_n9821_ ^ new_n6973_;
  assign n1257 = new_n6903_ | new_n6796_;
  assign new_n9801_ = ~new_n9986_ ^ new_n6974_;
  assign n1252 = new_n6904_ | new_n6797_;
  assign new_n9810_ = new_n6341_ & new_n9813_;
  assign new_n9813_ = new_n7423_ | new_n6798_;
  assign new_n9815_ = new_n7203_ | new_n6799_;
  assign new_n7106_ = ~new_n8307_;
  assign n1247 = new_n6905_ | new_n6800_;
  assign new_n9834_ = ~new_n9835_ ^ new_n9836_;
  assign new_n9836_ = ~new_n7359_ ^ new_n7373_;
  assign n1242 = new_n6906_ | new_n6801_;
  assign new_n9849_ = new_n9850_ ^ new_n9851_;
  assign new_n9850_ = ~new_n9852_ ^ new_n9853_;
  assign n1237 = new_n6907_ | new_n6802_;
  assign new_n9864_ = ~new_n9865_ ^ new_n9866_;
  assign new_n9866_ = new_n9867_ ^ new_n7384_;
  assign n1232 = new_n6908_ | new_n6803_;
  assign new_n7107_ = ~new_n8397_;
  assign n1227 = new_n6909_ | new_n6804_;
  assign new_n9886_ = ~new_n9745_ ^ new_n6975_;
  assign n1222 = new_n6910_ | new_n6805_;
  assign new_n9897_ = new_n9898_ & new_n6590_;
  assign new_n9900_ = new_n6342_ & new_n7416_;
  assign new_n9898_ = new_n6911_ | new_n6806_;
  assign n1217 = new_n6912_ | new_n6807_;
  assign new_n9923_ = new_n9924_ ^ new_n9925_;
  assign new_n9924_ = new_n9926_ ^ new_n7383_;
  assign n1212 = new_n6913_ | new_n6808_;
  assign new_n9296_ = new_n10319_ & new_n7264_;
  assign new_n9940_ = new_n9909_ | new_n7441_;
  assign new_n9943_ = new_n9945_ & new_n7441_;
  assign new_n9946_ = new_n7441_ ^ new_n9945_;
  assign n1207 = new_n6914_ | new_n6809_;
  assign new_n9957_ = ~new_n6951_ ^ new_n7346_;
  assign new_n9726_ = new_n7555_ | n1332;
  assign n1202 = new_n6915_ | new_n6810_;
  assign new_n9968_ = new_n9969_ ^ new_n9970_;
  assign new_n9969_ = ~new_n7220_ ^ new_n7375_;
  assign n1197 = new_n6916_ | new_n6811_;
  assign new_n7108_ = ~new_n9296_;
  assign new_n9983_ = ~new_n9567_ ^ new_n6976_;
  assign n1192 = new_n6917_ | new_n6812_;
  assign new_n9997_ = new_n9998_ & new_n6598_;
  assign new_n9694_ = new_n7299_ & new_n6599_;
  assign new_n9998_ = new_n7204_ | new_n6813_;
  assign new_n10004_ = ~new_n7315_ ^ new_n7569_;
  assign new_n10007_ = ~new_n9685_ ^ new_n7315_;
  assign new_n10014_ = new_n7373_ | new_n7359_;
  assign new_n9835_ = new_n6959_ ^ new_n7569_;
  assign new_n10022_ = new_n7374_ | new_n7360_;
  assign new_n8942_ = new_n10511_ & new_n10389_;
  assign new_n9609_ = new_n6960_ ^ new_n7569_;
  assign new_n10030_ = new_n7383_ | new_n9925_;
  assign new_n9926_ = new_n6343_ & new_n7153_;
  assign new_n10032_ = ~new_n7316_ ^ new_n7569_;
  assign new_n10035_ = ~new_n9685_ ^ new_n7316_;
  assign new_n9740_ = new_n7295_ & new_n6600_;
  assign new_n10041_ = ~new_n7319_ ^ new_n7569_;
  assign new_n10044_ = new_n9660_ | new_n9661_;
  assign new_n9661_ = new_n10049_ & new_n6602_;
  assign new_n10053_ = ~new_n7317_ ^ new_n7569_;
  assign new_n7109_ = ~new_n8942_;
  assign new_n10056_ = ~new_n9685_ ^ new_n7317_;
  assign new_n9817_ = new_n7300_ & new_n6603_;
  assign new_n10062_ = ~new_n7318_ ^ new_n7569_;
  assign new_n10065_ = new_n7378_ | new_n10069_;
  assign new_n10071_ = ~new_n9685_ ^ new_n7318_;
  assign new_n10049_ = new_n7375_ | new_n9970_;
  assign new_n9970_ = new_n6961_ ^ new_n7569_;
  assign new_n9660_ = new_n6962_ ^ new_n7569_;
  assign new_n10084_ = ~new_n9685_ ^ new_n7319_;
  assign new_n9925_ = new_n6963_ ^ new_n7569_;
  assign new_n7110_ = ~new_n10482_;
  assign new_n10094_ = ~new_n7320_ ^ new_n7569_;
  assign new_n10097_ = ~new_n9685_ ^ new_n7320_;
  assign n1187 = new_n6918_ | new_n6814_;
  assign new_n9547_ = new_n6344_ & new_n10109_;
  assign new_n9548_ = new_n6345_ & new_n10109_;
  assign new_n10114_ = new_n6346_ & new_n10122_;
  assign new_n10116_ = new_n6919_ | new_n6815_;
  assign new_n10127_ = new_n7187_ & new_n10703_;
  assign new_n10137_ = new_n7418_ & new_n7547_;
  assign new_n10126_ = new_n10139_ ^ new_n10069_;
  assign new_n9842_ = REG3_REG_4_ & n1332;
  assign new_n10069_ = new_n6964_ ^ new_n7569_;
  assign new_n10139_ = ~new_n7221_ ^ new_n7378_;
  assign new_n10149_ = ~new_n7328_ ^ new_n7569_;
  assign new_n10156_ = ~new_n7329_ ^ new_n7569_;
  assign new_n10155_ = new_n7188_ & new_n7169_;
  assign new_n10163_ = ~new_n7327_ ^ new_n7569_;
  assign new_n9867_ = new_n7161_ & new_n6606_;
  assign new_n10171_ = new_n7312_ | new_n7099_;
  assign new_n10178_ = new_n9851_ | new_n9852_;
  assign new_n9852_ = new_n6347_ & new_n7154_;
  assign new_n7034_ = ~new_n8247_;
  assign new_n7111_ = ~new_n9842_;
  assign new_n10184_ = ~new_n7321_ ^ new_n7569_;
  assign new_n10187_ = ~new_n9685_ ^ new_n7321_;
  assign new_n9640_ = new_n7301_ & new_n6609_;
  assign new_n10194_ = ~new_n7322_ ^ new_n7569_;
  assign new_n10199_ = new_n7377_ | new_n10201_;
  assign new_n10202_ = ~new_n9685_ ^ new_n7322_;
  assign new_n10207_ = ~new_n7323_ ^ new_n7569_;
  assign new_n10210_ = ~new_n9685_ ^ new_n7323_;
  assign new_n9851_ = new_n6965_ ^ new_n7569_;
  assign new_n10177_ = new_n9803_ & new_n10172_;
  assign new_n7112_ = ~new_n11060_;
  assign new_n10218_ = ~new_n7324_ ^ new_n7569_;
  assign new_n9803_ = new_n7175_ | new_n10173_;
  assign new_n10173_ = new_n6966_ ^ new_n7569_;
  assign new_n10227_ = ~new_n9685_ ^ new_n7325_;
  assign new_n10230_ = ~new_n9685_ ^ new_n7324_;
  assign new_n10235_ = ~new_n7325_ ^ new_n7569_;
  assign new_n10240_ = ~new_n7326_ ^ new_n7569_;
  assign new_n10243_ = ~new_n9685_ ^ new_n7326_;
  assign new_n10166_ = new_n7384_ | new_n9865_;
  assign new_n9865_ = new_n6967_ ^ new_n7569_;
  assign new_n7113_ = ~new_n8899_;
  assign new_n10253_ = ~new_n9685_ ^ new_n7327_;
  assign new_n9909_ = new_n7400_ | new_n9945_;
  assign new_n9945_ = new_n6968_ ^ new_n7569_;
  assign new_n10152_ = new_n7416_ & new_n7306_;
  assign new_n10263_ = ~new_n9685_ ^ new_n7328_;
  assign new_n10268_ = ~new_n9685_ ^ new_n7329_;
  assign new_n10145_ = new_n7376_ | new_n9595_;
  assign new_n9595_ = new_n6969_ ^ new_n7569_;
  assign new_n10277_ = new_n10703_ & new_n9269_;
  assign new_n10281_ = new_n6920_ | new_n7215_;
  assign new_n7114_ = ~new_n8989_;
  assign new_n10291_ = D_REG_29_ | D_REG_2_;
  assign new_n10290_ = D_REG_30_ | D_REG_31_;
  assign new_n10292_ = D_REG_23_ | D_REG_24_;
  assign new_n10297_ = D_REG_3_ | D_REG_4_;
  assign new_n10296_ = D_REG_5_ | D_REG_6_;
  assign new_n10299_ = D_REG_18_ | D_REG_19_;
  assign new_n10298_ = D_REG_20_ | D_REG_21_;
  assign new_n10306_ = D_REG_14_ | D_REG_15_;
  assign new_n10305_ = D_REG_16_ | D_REG_17_;
  assign new_n10308_ = D_REG_10_ | D_REG_11_;
  assign new_n10109_ = new_n10702_ & new_n10135_;
  assign new_n10307_ = D_REG_12_ | D_REG_13_;
  assign new_n10313_ = D_REG_28_ | D_REG_7_;
  assign new_n10312_ = D_REG_8_ | D_REG_9_;
  assign new_n10314_ = D_REG_26_ | D_REG_27_;
  assign new_n10315_ = new_n7410_ | D_REG_1_;
  assign new_n10317_ = new_n7410_ | D_REG_0_;
  assign new_n8432_ = ~B_REG;
  assign new_n10322_ = new_n7264_ & new_n7269_;
  assign n1182 = ~new_n6170_ | ~new_n5896_;
  assign new_n8450_ = new_n7118_ & new_n7701_;
  assign new_n7115_ = ~new_n10109_;
  assign new_n10332_ = new_n7550_ & new_n6612_;
  assign new_n10370_ = new_n6921_ | new_n6816_;
  assign new_n10374_ = new_n7529_ & new_n7485_;
  assign new_n10381_ = new_n7485_ & new_n10382_;
  assign new_n10382_ = new_n10383_ & new_n7529_;
  assign new_n10388_ = new_n10390_ & new_n6613_;
  assign new_n10397_ = new_n6922_ | new_n6817_;
  assign new_n10401_ = new_n7216_ | new_n6818_;
  assign new_n10369_ = new_n7515_ & new_n7542_;
  assign new_n10367_ = new_n7452_ & new_n7541_;
  assign new_n8890_ = new_n7248_ & new_n7445_;
  assign new_n10365_ = new_n7523_ & new_n7478_;
  assign new_n10363_ = new_n7409_ & new_n7406_;
  assign new_n10359_ = new_n7408_ & new_n7484_;
  assign new_n10357_ = new_n7479_ & new_n7546_;
  assign new_n10355_ = new_n7530_ & new_n7526_;
  assign new_n10350_ = new_n7422_ & new_n7477_;
  assign new_n10348_ = new_n7487_ & new_n7543_;
  assign new_n10346_ = new_n7514_ & new_n7413_;
  assign new_n10344_ = new_n7462_ & new_n7539_;
  assign new_n10340_ = new_n10420_ & new_n10421_;
  assign new_n7116_ = ~new_n8890_;
  assign new_n10422_ = ~new_n6952_ ^ new_n7701_;
  assign new_n8650_ = new_n7474_ & new_n7530_;
  assign new_n8564_ = new_n7477_ & new_n7487_;
  assign new_n8584_ = new_n7522_ & new_n7422_;
  assign new_n8742_ = new_n7486_ & new_n7484_;
  assign new_n8762_ = new_n7406_ & new_n7307_;
  assign new_n8710_ = new_n7408_ & new_n7479_;
  assign new_n10441_ = new_n7427_ & new_n10421_;
  assign new_n8532_ = new_n7543_ & new_n7514_;
  assign new_n8467_ = new_n7539_ & new_n7524_;
  assign new_n8980_ = new_n7251_ & new_n7393_;
  assign new_n9089_ = new_n7403_ & new_n7471_;
  assign new_n10454_ = new_n9228_ | new_n7411_;
  assign new_n9228_ = ~new_n9240_;
  assign new_n9240_ = ~new_n8257_ ^ new_n9216_;
  assign new_n9208_ = new_n7476_ & new_n10405_;
  assign new_n8880_ = new_n7515_ & new_n7470_;
  assign new_n8911_ = new_n7302_ & new_n7529_;
  assign new_n8853_ = new_n7542_ & new_n7541_;
  assign new_n10461_ = new_n8789_ & new_n8824_;
  assign new_n10463_ = new_n7428_ | new_n7275_;
  assign new_n7117_ = ~new_n8980_;
  assign new_n8940_ = new_n7485_ & new_n7289_;
  assign new_n10468_ = new_n7314_ | new_n10470_;
  assign new_n10470_ = new_n6923_ | new_n6819_;
  assign new_n8621_ = new_n7259_ & new_n7474_;
  assign new_n10496_ = new_n7486_ | new_n10416_;
  assign new_n10489_ = new_n6348_ & new_n7422_;
  assign new_n8586_ = new_n8627_ & new_n10495_;
  assign new_n8627_ = new_n10498_ & new_n7484_;
  assign new_n10498_ = new_n7408_ & new_n7365_;
  assign new_n10504_ = new_n7478_ & new_n7542_;
  assign new_n7035_ = ~new_n8265_;
  assign new_n10130_ = new_n11129_ | new_n9278_;
  assign new_n10501_ = new_n6924_ | new_n6820_;
  assign new_n8910_ = new_n6349_ & new_n7289_;
  assign new_n10389_ = new_n7453_ & new_n7415_;
  assign new_n10511_ = new_n7366_ & new_n7458_;
  assign new_n9090_ = new_n7472_ & new_n6614_;
  assign new_n10516_ = new_n7525_ | new_n9122_;
  assign new_n10515_ = new_n7520_ & new_n7473_;
  assign new_n10390_ = new_n7417_ & new_n7403_;
  assign new_n9184_ = new_n6350_ & new_n10405_;
  assign new_n9207_ = new_n7216_ & new_n7414_;
  assign new_n7118_ = ~new_n10130_;
  assign new_n9227_ = new_n10522_ & new_n6616_;
  assign new_n10522_ = new_n7506_ | new_n7549_;
  assign new_n10510_ = new_n7485_ & new_n7198_;
  assign new_n10383_ = new_n7475_ | new_n8968_;
  assign new_n10527_ = new_n10420_ & new_n7469_;
  assign new_n10539_ = new_n6925_ | new_n6821_;
  assign new_n10553_ = new_n7414_ & new_n8274_;
  assign new_n10405_ = new_n8262_ | new_n7531_;
  assign new_n10544_ = new_n6351_ & new_n7415_;
  assign new_n10556_ = new_n6352_ & new_n7417_;
  assign new_n7119_ = ~new_n7725_;
  assign new_n10538_ = new_n6928_ | new_n6822_;
  assign new_n10563_ = new_n6927_ | new_n6823_;
  assign new_n10566_ = new_n6926_ | new_n6824_;
  assign new_n10584_ = new_n6353_ & new_n7474_;
  assign new_n10589_ = new_n10635_ | DATAI_1_;
  assign new_n10592_ = new_n10635_ | DATAI_4_;
  assign new_n10590_ = new_n7476_ & new_n7414_;
  assign new_n10595_ = new_n10635_ | DATAI_2_;
  assign new_n10598_ = new_n10635_ | DATAI_3_;
  assign new_n10601_ = new_n7303_ & new_n7208_;
  assign new_n7120_ = ~new_n7728_;
  assign new_n10608_ = new_n10635_ | DATAI_5_;
  assign new_n10610_ = new_n10635_ | DATAI_8_;
  assign new_n10613_ = new_n10635_ | DATAI_7_;
  assign new_n10616_ = new_n10635_ | DATAI_9_;
  assign new_n10619_ = new_n10635_ | DATAI_6_;
  assign new_n10604_ = new_n10384_ & new_n7155_;
  assign new_n10625_ = new_n7487_ | new_n8502_;
  assign new_n10420_ = new_n7815_ | new_n7461_;
  assign new_n10421_ = new_n7480_ | new_n7407_;
  assign new_n10334_ = new_n7521_ | new_n7431_;
  assign new_n7731_ = new_n7739_ & new_n7738_;
  assign new_n10342_ = new_n7392_ & new_n7524_;
  assign new_n10633_ = new_n7208_ & new_n6617_;
  assign new_n10352_ = new_n7482_ & new_n7522_;
  assign new_n10495_ = new_n10643_ & new_n7530_;
  assign new_n10643_ = new_n7482_ & new_n7526_;
  assign new_n10648_ = new_n10635_ | DATAI_10_;
  assign new_n10651_ = new_n10635_ | DATAI_11_;
  assign new_n10657_ = new_n10635_ | DATAI_15_;
  assign new_n10659_ = IR_REG_15_ | IR_REG_31_;
  assign new_n10662_ = new_n10635_ | DATAI_16_;
  assign new_n7121_ = ~new_n7731_;
  assign new_n10667_ = new_n9417_ & IR_REG_16_;
  assign new_n10670_ = new_n10635_ | DATAI_12_;
  assign new_n10668_ = new_n7523_ & new_n7529_;
  assign new_n10672_ = new_n10635_ | DATAI_13_;
  assign new_n10674_ = IR_REG_13_ | IR_REG_31_;
  assign new_n10677_ = new_n10635_ | DATAI_17_;
  assign new_n10679_ = IR_REG_17_ | IR_REG_31_;
  assign new_n10680_ = new_n7528_ | new_n9410_;
  assign new_n9410_ = IR_REG_17_ & new_n7309_;
  assign new_n10361_ = new_n7486_ & new_n7307_;
  assign new_n7122_ = ~new_n8418_;
  assign new_n10684_ = new_n10635_ | DATAI_18_;
  assign new_n10691_ = new_n10635_ | DATAI_19_;
  assign new_n10693_ = new_n10635_ | DATAI_14_;
  assign new_n10697_ = new_n9432_ & IR_REG_14_;
  assign new_n10698_ = new_n6354_ & new_n10700_;
  assign new_n10700_ = new_n7115_ | new_n6825_;
  assign new_n10702_ = new_n9278_ & new_n10703_;
  assign n1178 = ~new_n6171_ | ~new_n5933_;
  assign n1174 = ~new_n6172_ | ~new_n5934_;
  assign n1170 = ~new_n6173_ | ~new_n5935_;
  assign new_n8895_ = new_n8083_ & new_n8928_;
  assign new_n7815_ = new_n6929_ | new_n6826_;
  assign new_n7797_ = new_n10730_ & REG3_REG_28_;
  assign new_n10730_ = new_n10740_ & REG3_REG_27_;
  assign n1166 = ~new_n6174_ | ~new_n5936_;
  assign new_n7816_ = ~new_n6953_ ^ REG3_REG_28_;
  assign n1162 = ~new_n6175_ | ~new_n5937_;
  assign new_n7833_ = ~new_n7338_ ^ REG3_REG_27_;
  assign n1158 = ~new_n6176_ | ~new_n5938_;
  assign new_n7850_ = new_n6355_ & new_n7338_;
  assign new_n10758_ = new_n10761_ & REG3_REG_25_;
  assign new_n7123_ = ~new_n8895_;
  assign new_n10759_ = ~REG3_REG_26_;
  assign n1154 = ~new_n6177_ | ~new_n5939_;
  assign new_n7867_ = ~new_n7339_ ^ REG3_REG_25_;
  assign n1150 = ~new_n6178_ | ~new_n5940_;
  assign new_n7884_ = new_n6356_ & new_n7339_;
  assign new_n10779_ = new_n7439_ & REG3_REG_23_;
  assign new_n10781_ = ~REG3_REG_24_;
  assign n1146 = ~new_n6179_ | ~new_n5941_;
  assign new_n7901_ = new_n7439_ ^ REG3_REG_23_;
  assign n1142 = ~new_n6180_ | ~new_n5942_;
  assign new_n8985_ = new_n8136_ & new_n9025_;
  assign new_n10799_ = new_n10800_ & new_n7213_;
  assign new_n10800_ = ~REG3_REG_22_;
  assign n1138 = ~new_n6181_ | ~new_n5943_;
  assign new_n7935_ = REG3_REG_21_ ^ new_n10810_;
  assign n1134 = ~new_n6182_ | ~new_n5944_;
  assign new_n7952_ = new_n6357_ & new_n7092_;
  assign new_n10820_ = new_n10822_ & REG3_REG_19_;
  assign new_n10821_ = ~REG3_REG_20_;
  assign n1130 = ~new_n6183_ | ~new_n5945_;
  assign new_n7969_ = ~REG3_REG_19_ ^ new_n7355_;
  assign new_n7036_ = ~new_n8281_;
  assign new_n7124_ = ~new_n8985_;
  assign n1126 = ~new_n6184_ | ~new_n5946_;
  assign new_n7986_ = new_n6358_ & new_n7355_;
  assign new_n10840_ = REG3_REG_18_ & REG3_REG_17_;
  assign new_n10841_ = ~REG3_REG_18_;
  assign n1122 = ~new_n6185_ | ~new_n5947_;
  assign new_n8003_ = ~new_n7340_ ^ REG3_REG_17_;
  assign n1118 = ~new_n6186_ | ~new_n5948_;
  assign new_n8020_ = new_n6359_ & new_n7340_;
  assign new_n10861_ = REG3_REG_16_ & REG3_REG_15_;
  assign new_n10863_ = ~REG3_REG_16_;
  assign new_n8982_ = new_n7249_ & new_n7380_;
  assign n1114 = ~new_n6187_ | ~new_n5949_;
  assign new_n8037_ = REG3_REG_15_ ^ new_n7440_;
  assign n1110 = ~new_n6188_ | ~new_n5950_;
  assign new_n10884_ = new_n10882_ & REG3_REG_13_;
  assign n1106 = ~new_n6189_ | ~new_n5951_;
  assign new_n8071_ = ~new_n7430_ ^ REG3_REG_13_;
  assign n1102 = ~new_n6190_ | ~new_n5952_;
  assign new_n8088_ = new_n6360_ & new_n7430_;
  assign new_n10902_ = new_n10905_ & REG3_REG_11_;
  assign new_n10903_ = ~REG3_REG_12_;
  assign new_n7125_ = ~new_n8982_;
  assign n1098 = ~new_n6191_ | ~new_n5953_;
  assign new_n8105_ = ~new_n7341_ ^ REG3_REG_11_;
  assign n1094 = ~new_n6192_ | ~new_n5954_;
  assign new_n8124_ = new_n6361_ & new_n7341_;
  assign new_n10923_ = new_n10926_ & REG3_REG_10_;
  assign new_n10924_ = ~REG3_REG_10_;
  assign n1090 = ~new_n6193_ | ~new_n5955_;
  assign new_n8141_ = ~new_n7342_ ^ REG3_REG_9_;
  assign n1086 = ~new_n6194_ | ~new_n5956_;
  assign new_n8159_ = new_n6362_ & new_n7342_;
  assign new_n7126_ = ~new_n9239_;
  assign new_n10944_ = new_n10945_ & REG3_REG_7_;
  assign new_n10946_ = ~REG3_REG_8_;
  assign n1082 = ~new_n6195_ | ~new_n5957_;
  assign new_n8176_ = new_n10945_ ^ REG3_REG_7_;
  assign new_n10945_ = new_n10956_ & REG3_REG_6_;
  assign new_n10956_ = new_n10966_ & REG3_REG_5_;
  assign n1078 = ~new_n6196_ | ~new_n5958_;
  assign new_n8194_ = ~new_n6954_ ^ REG3_REG_6_;
  assign n1074 = ~new_n6197_ | ~new_n5959_;
  assign new_n8211_ = ~new_n7343_ ^ REG3_REG_5_;
  assign new_n7594_ = REG3_REG_14_ & n1332;
  assign n1070 = ~new_n6198_ | ~new_n5960_;
  assign new_n8222_ = new_n10983_ & new_n7343_;
  assign new_n10983_ = REG3_REG_4_ | REG3_REG_3_;
  assign n1066 = ~new_n6199_ | ~new_n5961_;
  assign new_n8262_ = new_n6930_ | new_n6827_;
  assign new_n8244_ = ~REG3_REG_3_;
  assign n1062 = ~new_n6200_ | ~new_n5962_;
  assign n1058 = ~new_n6201_ | ~new_n5963_;
  assign n1054 = ~new_n6202_ | ~new_n5964_;
  assign n1050 = new_n6931_ | new_n6828_;
  assign new_n7127_ = ~new_n7594_;
  assign new_n11015_ = new_n7206_ | new_n7100_;
  assign new_n11014_ = new_n11018_ & new_n11019_;
  assign new_n11019_ = new_n7548_ | new_n6829_;
  assign new_n11021_ = REG1_REG_0_ | IR_REG_0_;
  assign new_n11018_ = new_n7488_ | new_n6830_;
  assign n1046 = new_n6932_ | new_n6831_;
  assign new_n11029_ = new_n7554_ | new_n11036_;
  assign new_n11032_ = ~new_n7364_ ^ new_n11034_;
  assign new_n11034_ = ~new_n11035_ ^ new_n7426_;
  assign new_n11037_ = ~new_n7432_ ^ new_n11038_;
  assign new_n7697_ = REG3_REG_19_ & n1332;
  assign new_n11038_ = ~new_n11039_ ^ new_n7426_;
  assign n1042 = new_n6933_ | new_n6832_;
  assign new_n11049_ = ~new_n11050_ ^ new_n11341_;
  assign new_n11051_ = ~new_n11052_ ^ new_n11417_;
  assign new_n11056_ = ~REG1_REG_2_ ^ new_n11417_;
  assign new_n11054_ = new_n6363_ & new_n7554_;
  assign new_n11058_ = ~new_n11341_ ^ REG2_REG_2_;
  assign n1038 = new_n6934_ | new_n6833_;
  assign new_n11068_ = new_n6364_ & new_n7554_;
  assign new_n11072_ = ~new_n7504_ ^ new_n11074_;
  assign new_n7128_ = ~new_n7697_;
  assign new_n11077_ = new_n7548_ | new_n7192_;
  assign new_n11080_ = ~REG2_REG_3_ ^ new_n7504_;
  assign n1034 = new_n6935_ | new_n6834_;
  assign new_n11089_ = ~REG1_REG_4_ ^ new_n7349_;
  assign new_n11087_ = new_n6365_ & new_n7554_;
  assign new_n11092_ = ~new_n7503_ ^ new_n11094_;
  assign new_n11098_ = ~REG2_REG_4_ ^ new_n7503_;
  assign new_n11099_ = ~new_n11090_ ^ REG1_REG_4_;
  assign new_n11105_ = new_n7390_ | REG2_REG_0_;
  assign new_n11104_ = new_n11107_ & new_n6624_;
  assign new_n7632_ = REG3_REG_16_ & n1332;
  assign new_n11107_ = new_n9873_ | new_n11106_;
  assign new_n9873_ = new_n10201_ ^ new_n11109_;
  assign new_n11109_ = ~new_n9685_ ^ new_n7377_;
  assign new_n10201_ = new_n6970_ ^ new_n7569_;
  assign new_n9272_ = new_n7263_ & new_n7314_;
  assign new_n9292_ = new_n11129_ & new_n7550_;
  assign new_n11130_ = new_n10635_ | DATAI_0_;
  assign new_n10709_ = new_n11137_ & new_n7424_;
  assign new_n11137_ = ~new_n11138_;
  assign new_n10729_ = new_n7424_ & new_n11138_;
  assign new_n7129_ = ~new_n7632_;
  assign new_n11138_ = ~IR_REG_30_ ^ new_n9536_;
  assign new_n9681_ = new_n6366_ & new_n7451_;
  assign new_n11151_ = IR_REG_19_ | IR_REG_31_;
  assign new_n11152_ = new_n7527_ | new_n9396_;
  assign new_n9396_ = IR_REG_19_ & new_n7308_;
  assign new_n11153_ = STATE_REG & new_n7450_;
  assign n1030 = new_n6936_ | new_n6835_;
  assign new_n11161_ = new_n6367_ & new_n7554_;
  assign new_n11165_ = ~new_n7494_ ^ new_n11167_;
  assign new_n11170_ = new_n7548_ | new_n7193_;
  assign new_n7037_ = ~new_n9948_;
  assign new_n7653_ = REG3_REG_17_ & n1332;
  assign new_n11173_ = ~REG2_REG_5_ ^ new_n7494_;
  assign n1026 = new_n6937_ | new_n6836_;
  assign new_n11183_ = ~REG1_REG_6_ ^ new_n7499_;
  assign new_n11181_ = new_n6368_ & new_n7554_;
  assign new_n11186_ = ~new_n7502_ ^ new_n11188_;
  assign new_n11192_ = ~REG2_REG_6_ ^ new_n7502_;
  assign new_n11193_ = ~new_n7499_ ^ new_n11194_;
  assign n1022 = new_n6938_ | new_n6837_;
  assign new_n11203_ = ~REG2_REG_7_ ^ new_n7498_;
  assign new_n11205_ = ~new_n11206_ ^ new_n11381_;
  assign new_n7130_ = ~new_n7653_;
  assign new_n11210_ = ~new_n11381_ ^ REG1_REG_7_;
  assign new_n11208_ = new_n6369_ & new_n7554_;
  assign new_n11212_ = ~new_n7498_ ^ new_n11213_;
  assign n1018 = new_n6939_ | new_n6838_;
  assign new_n11220_ = new_n6370_ & new_n7554_;
  assign new_n11224_ = ~new_n7501_ ^ new_n11226_;
  assign new_n11229_ = new_n7548_ | new_n7194_;
  assign new_n11232_ = ~REG2_REG_8_ ^ new_n7501_;
  assign n1014 = new_n6940_ | new_n6839_;
  assign new_n11241_ = ~REG2_REG_9_ ^ new_n7497_;
  assign new_n7572_ = REG3_REG_13_ & n1332;
  assign new_n11243_ = ~new_n11248_ ^ REG1_REG_9_;
  assign new_n11247_ = ~REG1_REG_9_ ^ new_n7348_;
  assign new_n11245_ = new_n6371_ & new_n7554_;
  assign new_n11250_ = ~new_n7497_ ^ new_n11251_;
  assign n1010 = new_n6941_ | new_n6840_;
  assign new_n11258_ = new_n6372_ & new_n7554_;
  assign new_n11262_ = ~new_n7500_ ^ new_n11264_;
  assign new_n11267_ = new_n7548_ | new_n7195_;
  assign new_n11270_ = ~REG2_REG_10_ ^ new_n7500_;
  assign n1006 = new_n6942_ | new_n6841_;
  assign new_n7131_ = ~new_n7572_;
  assign new_n11279_ = ~REG2_REG_11_ ^ new_n7496_;
  assign new_n11281_ = ~new_n7495_ ^ new_n11283_;
  assign new_n11287_ = ~REG1_REG_11_ ^ new_n7495_;
  assign new_n11285_ = new_n6373_ & new_n7554_;
  assign new_n11289_ = ~new_n7496_ ^ new_n11290_;
  assign n1002 = new_n6943_ | new_n6842_;
  assign new_n11300_ = ~new_n7738_ ^ REG1_REG_12_;
  assign new_n11298_ = new_n6374_ & new_n7554_;
  assign new_n11302_ = ~new_n7505_ ^ new_n7766_;
  assign new_n7766_ = ~REG2_REG_12_;
  assign new_n7675_ = REG3_REG_18_ & n1332;
  assign new_n11307_ = new_n9447_ & IR_REG_12_;
  assign new_n11310_ = ~REG2_REG_12_ ^ new_n7505_;
  assign new_n11290_ = ~REG2_REG_11_;
  assign new_n11313_ = new_n7496_ | new_n7460_;
  assign new_n11264_ = ~REG2_REG_10_;
  assign new_n11316_ = new_n7500_ | new_n7448_;
  assign new_n11251_ = ~REG2_REG_9_;
  assign new_n11319_ = new_n7497_ | new_n7516_;
  assign new_n11226_ = ~REG2_REG_8_;
  assign new_n11322_ = new_n7501_ | new_n7449_;
  assign new_n7132_ = ~new_n7675_;
  assign new_n11213_ = ~REG2_REG_7_;
  assign new_n11325_ = new_n7498_ | new_n7517_;
  assign new_n11188_ = ~REG2_REG_6_;
  assign new_n11328_ = new_n7502_ | new_n11179_;
  assign new_n11167_ = ~REG2_REG_5_;
  assign new_n11331_ = new_n7494_ | new_n11159_;
  assign new_n11094_ = ~REG2_REG_4_;
  assign new_n11334_ = new_n7503_ | new_n7511_;
  assign new_n11074_ = ~REG2_REG_3_;
  assign new_n11337_ = new_n7504_ | new_n11066_;
  assign new_n7613_ = REG3_REG_15_ & n1332;
  assign new_n11050_ = ~REG2_REG_2_;
  assign new_n11035_ = ~REG2_REG_1_;
  assign new_n11344_ = new_n7364_ | new_n11036_;
  assign new_n11345_ = new_n11017_ & new_n11106_;
  assign new_n11346_ = ~REG1_REG_12_ ^ new_n7350_;
  assign new_n11283_ = ~REG1_REG_11_;
  assign new_n11347_ = new_n7495_ | new_n10652_;
  assign new_n11351_ = IR_REG_11_ | IR_REG_31_;
  assign new_n11356_ = REG1_REG_9_ & new_n7209_;
  assign new_n11362_ = new_n7209_ & new_n6631_;
  assign new_n7133_ = ~new_n7613_;
  assign new_n11364_ = ~REG1_REG_9_;
  assign new_n11366_ = IR_REG_31_ | IR_REG_9_;
  assign new_n11370_ = new_n6375_ & new_n11373_;
  assign new_n11231_ = new_n11373_ | new_n6843_;
  assign new_n11206_ = ~REG1_REG_7_;
  assign new_n11194_ = ~REG1_REG_6_;
  assign new_n11382_ = new_n7499_ | new_n7402_;
  assign new_n11392_ = REG1_REG_4_ & new_n7210_;
  assign new_n9499_ = new_n6376_ & new_n9492_;
  assign new_n11398_ = new_n7210_ & new_n6633_;
  assign new_n9724_ = new_n10194_ & new_n10195_;
  assign new_n11400_ = ~REG1_REG_4_;
  assign new_n11406_ = new_n6377_ & new_n11409_;
  assign new_n9516_ = ~IR_REG_3_;
  assign new_n11079_ = new_n11409_ | new_n6844_;
  assign new_n11052_ = ~REG1_REG_2_;
  assign new_n11039_ = ~REG1_REG_1_;
  assign new_n11420_ = new_n11036_ | new_n7432_;
  assign new_n11409_ = ~REG1_REG_3_;
  assign new_n11373_ = ~REG1_REG_8_;
  assign new_n9537_ = new_n6378_ & STATE_REG;
  assign new_n7134_ = ~new_n9724_;
  assign new_n11439_ = IR_REG_21_ | IR_REG_31_;
  assign new_n9338_ = ~IR_REG_27_;
  assign new_n9329_ = ~IR_REG_28_;
  assign new_n11457_ = IR_REG_23_ | IR_REG_31_;
  assign n1332 = ~STATE_REG;
  assign new_n11464_ = new_n7401_ & IR_REG_25_;
  assign new_n11459_ = new_n7260_ & new_n10323_;
  assign new_n9536_ = ~IR_REG_31_;
  assign new_n11471_ = IR_REG_26_ & new_n7313_;
  assign new_n9351_ = ~IR_REG_25_;
  assign new_n7038_ = ~new_n9986_;
  assign new_n7135_ = ~new_n10546_;
  assign new_n9361_ = ~IR_REG_24_;
  assign new_n9376_ = ~IR_REG_22_;
  assign new_n9391_ = ~IR_REG_20_;
  assign new_n9405_ = ~IR_REG_18_;
  assign new_n9419_ = ~IR_REG_16_;
  assign new_n9434_ = ~IR_REG_14_;
  assign new_n9449_ = ~IR_REG_12_;
  assign new_n9464_ = ~IR_REG_10_;
  assign new_n9478_ = ~IR_REG_8_;
  assign new_n11431_ = ~IR_REG_7_;
  assign new_n9794_ = REG3_REG_5_ & n1332;
  assign new_n9494_ = ~IR_REG_6_;
  assign new_n9508_ = ~IR_REG_4_;
  assign new_n11427_ = ~IR_REG_2_;
  assign new_n9530_ = ~IR_REG_0_;
  assign new_n9532_ = ~IR_REG_1_;
  assign new_n10406_ = new_n7476_ & new_n5539_;
  assign new_n10399_ = new_n4935_ & new_n10401_;
  assign new_n10391_ = new_n4934_ & new_n7471_;
  assign new_n10385_ = new_n4936_ & new_n5538_;
  assign new_n10371_ = new_n4933_ & new_n7470_;
  assign new_n7136_ = ~new_n9794_;
  assign new_n10372_ = new_n10378_ & new_n5537_;
  assign new_n10558_ = new_n10525_ & new_n5566_;
  assign new_n10551_ = new_n7103_ & new_n5565_;
  assign new_n10572_ = new_n7470_ & new_n5569_;
  assign new_n10638_ = new_n4963_ & new_n7514_;
  assign new_n10630_ = new_n7539_ & new_n5575_;
  assign new_n10549_ = new_n10405_ & new_n5564_;
  assign new_n10546_ = new_n6384_ | new_n6423_;
  assign new_n10569_ = new_n10361_ & new_n5568_;
  assign new_n10603_ = new_n6386_ | new_n6424_;
  assign new_n9976_ = REG3_REG_6_ & n1332;
  assign new_n10628_ = new_n10420_ & new_n5574_;
  assign new_n10583_ = new_n10584_ & new_n5571_;
  assign new_n10554_ = new_n4949_ & new_n7475_;
  assign new_n10542_ = new_n4976_ & new_n5577_;
  assign new_n10565_ = new_n10566_ & new_n5567_;
  assign new_n10564_in = new_n4950_ & new_n7484_;
  assign new_n10640_ = new_n4964_ & new_n7522_;
  assign new_n10641_ = new_n10495_ & new_n5576_;
  assign new_n10602_ = new_n6385_ | new_n7214_;
  assign new_n10626_ = new_n10421_ & new_n5573_;
  assign new_n7137_in = ~new_n9976_;
  assign new_n10482_ = new_n8416_ & new_n5560_;
  assign new_n10540_ = new_n10384_ & new_n5563_;
  assign new_n10621_in = new_n4962_ & new_n5572_;
  assign new_n10487_in = new_n4945_ & new_n7487_;
  assign new_n11410_ = new_n7446_ & new_n6998_;
  assign new_n7725_in = new_n7605_ & new_n7057_;
  assign new_n8519_in = new_n4680_ & new_n7879_;
  assign new_n8670_in = new_n7456_ | new_n6418_;
  assign new_n9139_ = new_n4751_ & new_n9173_;
  assign new_n8628_ = new_n7233_ & new_n7896_;
  assign new_n9544_in = REG3_REG_7_ & n1332;
  assign new_n10229_ = new_n4915_ & new_n5516_;
  assign new_n10196_in = new_n4905_ & new_n5507_;
  assign new_n10186_ = new_n4902_ & new_n5503_;
  assign new_n10151_ = new_n4925_ & new_n5526_;
  assign new_n10034_in = new_n4874_ & new_n5475_;
  assign new_n10209_in = new_n4907_ & new_n5509_;
  assign new_n10055_ = new_n4878_ & new_n5478_;
  assign new_n10096_ = new_n4891_ & new_n5490_;
  assign new_n10006_in = new_n4866_ & new_n5466_;
  assign new_n9680_ = new_n6979_ & new_n7066_;
  assign new_n7138_ = ~new_n9544_;
  assign new_n10426_in = new_n4939_ & new_n5542_;
  assign new_n10536_ = new_n4951_ & new_n7469_;
  assign new_n10479_in = new_n6158_ & new_n5548_;
  assign new_n10471_ = new_n4944_ & new_n10334_;
  assign new_n11341_in = new_n5081_ & new_n5690_;
  assign new_n11415_ = new_n7149_ & new_n5701_;
  assign new_n11381_ = new_n11382_ & new_n5695_;
  assign new_n11374_ = new_n7517_ & new_n6997_;
  assign new_n7591_ = new_n4567_ & new_n7121_;
  assign new_n7728_ = new_n7576_ & new_n7062_;
  assign new_n9701_ = REG3_REG_8_ & n1332;
  assign new_n7610_ = new_n4573_ & new_n5134_;
  assign new_n7629_ = new_n4566_ & new_n7119_;
  assign new_n7628_ = REG1_REG_15_ & new_n5127_;
  assign new_n8671_in = new_n4696_ & new_n7152_;
  assign new_n8833_ = new_n4714_ & new_n6495_;
  assign new_n10413_ = new_n7381_ & new_n8805_;
  assign new_n8840_ = new_n7229_ & new_n7382_;
  assign new_n10452_ = new_n8154_ & new_n7251_;
  assign new_n10396_ = new_n7379_ & new_n9106_;
  assign new_n10393_ = new_n7236_ & new_n8189_;
  assign new_n7139_ = ~new_n9701_;
  assign new_n10404_ = new_n7238_ & new_n9172_;
  assign new_n9155_ = new_n7369_ & new_n9171_;
  assign new_n9242_ = new_n9243_ & new_n7065_;
  assign new_n10123_ = new_n9290_ & new_n6996_;
  assign new_n8440_ = new_n4669_ & new_n7539_;
  assign new_n8445_ = new_n4670_ & new_n7524_;
  assign new_n8443_ = new_n8454_ & new_n7519_;
  assign new_n8442_ = new_n7231_ & new_n7808_;
  assign new_n8473_ = new_n7845_ & new_n7239_;
  assign new_n8535_ = new_n7862_ & new_n7240_;
  assign new_n9857_ = REG3_REG_9_ & n1332;
  assign new_n10493_ = new_n8621_ & new_n5551_;
  assign new_n10433_ = new_n7879_ & new_n7391_;
  assign new_n8619_ = new_n8625_ & new_n5262_;
  assign new_n8613_ = new_n7474_ & new_n5260_;
  assign new_n8618_ = new_n7234_ & new_n7913_;
  assign new_n8623_ = new_n7930_ & new_n7241_;
  assign new_n10417_ = new_n8728_ & new_n7385_;
  assign new_n8711_ = new_n7438_ & new_n8729_;
  assign new_n8713_ = new_n7964_ & new_n7243_;
  assign new_n10414_ = new_n7370_ & new_n7998_;
  assign new_n9287_ = new_n10315_ & new_n7108_;
  assign new_n7140_ = ~new_n9857_;
  assign new_n10503_ = new_n10504_ & new_n5555_;
  assign new_n8777_ = new_n4709_ & new_n7101_;
  assign new_n8801_ = new_n4708_ & new_n5291_;
  assign new_n8820_ = new_n7532_ & new_n8841_;
  assign new_n8821_ = new_n8032_ & new_n7245_;
  assign new_n8857_ = new_n8049_ & new_n7229_;
  assign new_n10376_ = new_n7437_ & new_n8927_;
  assign new_n10460_ = new_n8066_ & new_n7246_;
  assign new_n8921_ = new_n4722_ & new_n8928_;
  assign new_n8924_ = new_n7180_ & new_n5311_;
  assign new_n9616_ = REG3_REG_10_ & n1332;
  assign new_n8941_ = new_n7458_ & new_n5559_;
  assign new_n8967_ = new_n7380_ & new_n9024_;
  assign new_n9005_ = new_n8136_ & new_n7250_;
  assign new_n9020_ = new_n7117_ & new_n5332_;
  assign new_n9091_ = new_n6383_ | new_n7151_;
  assign new_n9078_ = new_n7097_ & new_n5342_;
  assign new_n9102_ = new_n4745_ & new_n5341_;
  assign new_n9137_ = new_n4755_ & new_n7102_;
  assign new_n9167_ = new_n4754_ & new_n5351_;
  assign new_n10402_ = new_n9227_ & new_n7103_;
  assign new_n7141_ = ~new_n9616_;
  assign new_n10284_ = new_n4930_ & new_n5533_;
  assign new_n10283_ = new_n4931_ & new_n5534_;
  assign new_n9560_ = new_n10227_ & new_n6991_;
  assign new_n10154_ = new_n7158_ & new_n5499_;
  assign new_n10165_ = new_n4921_ & new_n5522_;
  assign new_n10242_ = new_n4917_ & new_n5518_;
  assign new_n9725_ = new_n10202_ & new_n6988_;
  assign new_n9741_ = new_n7071_ & new_n7153_;
  assign new_n10157_ = new_n4926_ & new_n5528_;
  assign new_n10064_ = new_n4880_ & new_n5481_;
  assign new_n9931_ = REG3_REG_11_ & n1332;
  assign new_n10221_ = new_n4909_ & new_n5511_;
  assign new_n10174_ = new_n4910_ & new_n5512_;
  assign new_n10118_ = new_n7450_ & new_n5494_;
  assign new_n9818_ = new_n7072_ & new_n7063_;
  assign new_n9647_ = new_n10187_ & new_n6987_;
  assign new_n11117_ = new_n5051_ & new_n7550_;
  assign new_n10132_ = new_n4895_ & new_n7547_;
  assign new_n10043_ = new_n4886_ & new_n5486_;
  assign new_n9902_ = new_n10263_ & new_n6994_;
  assign new_n9907_ = new_n4850_ & new_n7306_;
  assign new_n7142_ = ~new_n9931_;
  assign new_n9747_ = new_n10035_ & new_n6982_;
  assign new_n10260_ = new_n4923_ & new_n5524_;
  assign new_n9912_ = new_n7271_ & new_n5454_;
  assign new_n9645_ = new_n10210_ & new_n6989_;
  assign new_n9822_ = new_n10056_ & new_n6983_;
  assign new_n10220_ = new_n4913_ & new_n5514_;
  assign new_n9695_ = new_n10097_ & new_n6986_;
  assign new_n9776_ = new_n10007_ & new_n6981_;
  assign new_n10336_ = new_n7388_ & new_n5536_;
  assign new_n10337_ = new_n7521_ & new_n7431_;
  assign new_n9752_ = REG3_REG_12_ & n1332;
  assign new_n10446_ = new_n4942_ & new_n5544_;
  assign new_n10447_ = new_n4941_ & new_n5543_;
  assign new_n10427_ = new_n4938_ & new_n5541_;
  assign new_n10472_ = new_n4943_ & new_n5546_;
  assign new_n10134_ = new_n5052_ & new_n11129_;
  assign new_n11136_ = new_n5057_ & new_n5661_;
  assign new_n11073_ = new_n5080_ & new_n5689_;
  assign new_n11070_ = new_n7080_ & new_n11079_;
  assign new_n11093_ = new_n5079_ & new_n5688_;
  assign new_n11171_ = new_n5088_ & new_n7147_;
  assign new_n7143_ = ~new_n9752_;
  assign new_n11166_ = new_n5078_ & new_n5687_;
  assign new_n11187_ = new_n5077_ & new_n5686_;
  assign new_n11184_ = new_n7061_ & new_n5697_;
  assign new_n11204_ = new_n5076_ & new_n5685_;
  assign new_n11379_ = new_n7146_ & new_n5694_;
  assign new_n11225_ = new_n5075_ & new_n5684_;
  assign new_n11242_ = new_n5074_ & new_n5683_;
  assign new_n11268_ = new_n5083_ & new_n7144_;
  assign new_n11263_ = new_n5073_ & new_n5682_;
  assign new_n11280_ = new_n5072_ & new_n5681_;
  assign new_n11355_ = new_n10617_ & new_n7348_;
  assign new_n11282_ = new_n7060_ & new_n5692_;
  assign new_n7767_ = new_n5071_ & new_n5680_;
  assign new_n7587_ = new_n4574_ & new_n5135_;
  assign new_n7581_ = new_n7304_ & new_n7062_;
  assign new_n7626_ = new_n4572_ & new_n5133_;
  assign new_n7621_ = new_n7096_ & new_n7093_;
  assign new_n7643_ = new_n4571_ & new_n5132_;
  assign new_n7662_ = new_n4570_ & new_n5131_;
  assign new_n7664_ = new_n4565_ & new_n5125_;
  assign new_n7683_ = new_n4564_ & new_n5124_;
  assign new_n7144_ = ~new_n11355_;
  assign new_n7687_ = new_n4569_ & new_n5130_;
  assign new_n7706_ = new_n4568_ & new_n5129_;
  assign new_n7708_ = new_n4563_ & new_n5123_;
  assign new_n8456_ = new_n8481_ & new_n5236_;
  assign new_n8485_ = new_n4679_ & new_n5241_;
  assign new_n8549_ = new_n7177_ & new_n5247_;
  assign new_n8598_ = new_n8635_ & new_n5264_;
  assign new_n10780_ = new_n10800_ | new_n7213_;
  assign new_n8639_ = new_n8660_ & new_n5270_;
  assign new_n8660_ = new_n4692_ & new_n6478_;
  assign new_n11371_ = new_n11381_ & new_n10614_;
  assign new_n8835_ = new_n7282_ & new_n5302_;
  assign new_n10862_ = new_n7430_ | new_n6440_;
  assign new_n8867_ = new_n7058_ & new_n5307_;
  assign new_n8923_ = new_n7116_ & new_n5316_;
  assign new_n9018_ = new_n4734_ & new_n9025_;
  assign new_n9021_ = new_n7182_ & new_n5328_;
  assign new_n8255_ = new_n9234_ & new_n7442_;
  assign new_n11145_ = new_n5059_ & new_n6628_;
  assign new_n9196_ = new_n4761_ & new_n5359_;
  assign new_n10278_ = new_n9287_ & new_n7095_;
  assign new_n7039_ = ~new_n9287_;
  assign new_n7145_ = ~new_n11371_;
  assign new_n9274_ = new_n7069_ | new_n6420_;
  assign new_n8418_ = new_n4667_ & new_n5227_;
  assign new_n8478_ = new_n7808_ & new_n5235_;
  assign new_n8495_ = new_n4677_ & new_n5239_;
  assign new_n8471_ = new_n7477_ & new_n5244_;
  assign new_n8541_ = new_n7845_ & new_n5246_;
  assign new_n8585_ = new_n4946_ & new_n5550_;
  assign new_n8591_ = new_n7879_ & new_n5255_;
  assign new_n8609_ = new_n6380_ | new_n6417_;
  assign new_n8620_ = new_n8621_ & new_n5261_;
  assign new_n7146_ = ~new_n11374_;
  assign new_n8610_ = new_n8611_ & new_n5259_;
  assign new_n8617_ = new_n7546_ & new_n5267_;
  assign new_n8657_ = new_n7913_ & new_n5269_;
  assign new_n8709_ = new_n7486_ & new_n5276_;
  assign new_n8719_ = new_n7947_ & new_n5278_;
  assign new_n8714_ = new_n7307_ & new_n5552_;
  assign new_n8761_ = new_n7523_ & new_n5553_;
  assign new_n8767_ = new_n7981_ & new_n5286_;
  assign new_n8788_ = new_n10501_ & new_n5554_;
  assign new_n8817_ = new_n8824_ & new_n5294_;
  assign new_n11391_ = new_n10593_ & new_n7349_;
  assign new_n8830_ = new_n8015_ & new_n5296_;
  assign new_n8856_ = new_n7529_ & new_n5556_;
  assign new_n8885_ = new_n8049_ & new_n5306_;
  assign new_n8947_ = new_n8083_ & new_n5315_;
  assign new_n8964_ = new_n8971_ & new_n5319_;
  assign new_n8116_ = new_n8119_ & new_n5327_;
  assign new_n9006_ = new_n10512_ & new_n5557_;
  assign new_n10512_ = new_n4947_ & new_n6615_;
  assign new_n9036_ = new_n7415_ & new_n7475_;
  assign new_n9055_ = new_n4738_ & new_n7041_;
  assign new_n7147_ = ~new_n11391_;
  assign new_n8151_ = new_n8154_ & new_n5336_;
  assign new_n9060_ = new_n9090_ | new_n7197_;
  assign new_n9118_ = new_n4746_ & new_n7040_;
  assign new_n8186_ = new_n8189_ & new_n5346_;
  assign new_n9172_ = new_n4953_ & new_n10592_;
  assign new_n10523_ = new_n7389_ & new_n5558_;
  assign new_n8254_ = new_n8257_ & new_n5363_;
  assign new_n9256_ = new_n7288_ & new_n7065_;
  assign new_n9285_ = new_n6382_ | new_n6422_;
  assign new_n9255_ = new_n6980_ & new_n9235_;
  assign new_n11407_ = new_n11417_ & new_n10596_;
  assign new_n11441_ = new_n5097_ & new_n6636_;
  assign new_n9582_ = new_n4820_ & new_n7064_;
  assign new_n9583_ = new_n4821_ & new_n6578_;
  assign new_n9689_ = new_n4818_ & new_n5411_;
  assign new_n9596_ = new_n4899_ & new_n7274_;
  assign new_n10271_ = new_n4927_ & new_n5529_;
  assign new_n9597_ = new_n4928_ & new_n5530_;
  assign new_n10023_ = new_n4870_ & new_n5471_;
  assign new_n9612_ = new_n4872_ & new_n5472_;
  assign new_n9611_ = new_n4887_ & new_n5473_;
  assign new_n7148_ = ~new_n11407_;
  assign new_n9626_ = new_n10253_ & new_n6993_;
  assign new_n9641_ = new_n7074_ & new_n7154_;
  assign new_n9642_ = new_n4811_ & new_n7279_;
  assign new_n9662_ = new_n4875_ & new_n6601_;
  assign new_n10081_ = new_n4884_ & new_n5484_;
  assign new_n10050_ = new_n4881_ & new_n7220_;
  assign new_n9677_ = new_n4816_ & new_n5408_;
  assign new_n9676_ = new_n4817_ & new_n5409_;
  assign new_n9684_ = new_n4819_ & new_n5410_;
  assign new_n10170_ = new_n4911_ & new_n6607_;
  assign new_n7149_ = ~new_n11410_;
  assign new_n9712_ = new_n10243_ & new_n6992_;
  assign new_n9723_ = new_n4903_ & new_n5505_;
  assign new_n9742_ = new_n4828_ & new_n7278_;
  assign new_n9762_ = new_n10268_ & new_n5527_;
  assign new_n9789_ = new_n10071_ & new_n6984_;
  assign new_n9804_ = new_n10173_ & new_n7175_;
  assign new_n9819_ = new_n4838_ & new_n7273_;
  assign new_n9838_ = new_n4869_ & new_n5469_;
  assign new_n9837_ = new_n4871_ & new_n5470_;
  assign new_n10015_ = new_n4867_ & new_n5468_;
  assign new_n9343_ = new_n11471_ | new_n7481_;
  assign new_n9853_ = new_n4900_ & new_n6608_;
  assign new_n10215_ = new_n4908_ & new_n5510_;
  assign new_n10248_ = new_n4918_ & new_n5519_;
  assign new_n9868_ = new_n4919_ & new_n5520_;
  assign new_n10200_ = new_n11110_ & new_n5655_;
  assign new_n11110_ = new_n5049_ & new_n6625_;
  assign new_n11116_ = new_n5050_ & new_n6626_;
  assign new_n11115_ = new_n11120_ & new_n5656_;
  assign new_n11120_ = new_n5054_ & new_n6627_;
  assign new_n10121_ = new_n10128_ & new_n5495_;
  assign new_n7150_ = ~new_n9343_;
  assign new_n10128_ = new_n4896_ & new_n6605_;
  assign new_n9746_ = new_n10084_ & new_n6985_;
  assign new_n9899_ = new_n9900_ & new_n5446_;
  assign new_n9927_ = new_n4888_ & new_n5487_;
  assign new_n10091_ = new_n4889_ & new_n5488_;
  assign new_n9971_ = new_n4876_ & new_n7063_;
  assign new_n10076_ = new_n4882_ & new_n5482_;
  assign new_n9972_ = new_n4883_ & new_n5483_;
  assign new_n9563_ = new_n10230_ & new_n6990_;
  assign new_n10000_ = new_n7073_ & new_n7064_;
  assign new_n9156_ = new_n9184_ & new_n7459_;
  assign new_n10002_ = new_n4864_ & new_n7277_;
  assign new_n9568_ = new_n7798_ & new_n5531_;
  assign new_n10070_ = new_n4898_ & new_n5497_;
  assign new_n10068_ = new_n10145_ & new_n5498_;
  assign new_n10140_ = new_n4897_ & new_n5496_;
  assign new_n11446_ = new_n5098_ & new_n6637_;
  assign new_n11451_ = new_n5099_ & new_n6638_;
  assign new_n10333_ = new_n10334_ & new_n5535_;
  assign new_n10423_ = new_n4940_ & new_n5540_;
  assign new_n10466_ = new_n4948_ & new_n5561_;
  assign new_n7023_ = ~new_n8074_;
  assign new_n9120_ = new_n7473_ & new_n7472_;
  assign new_n7151_ = ~new_n9156_;
  assign new_n10467_ = new_n10468_ & new_n5545_;
  assign new_n10734_ = new_n4986_ & new_n5582_;
  assign new_n10733_ = new_n4987_ & new_n5583_;
  assign new_n10744_ = new_n4988_ & new_n5584_;
  assign new_n10743_ = new_n4989_ & new_n5585_;
  assign new_n10765_ = new_n4992_ & new_n5589_;
  assign new_n10764_ = new_n4993_ & new_n5590_;
  assign new_n10794_ = new_n4998_ & new_n5596_;
  assign new_n10793_ = new_n4999_ & new_n5597_;
  assign new_n10826_ = new_n5004_ & new_n5603_;
  assign new_n8696_ = new_n7947_ & new_n8728_;
  assign new_n10825_ = new_n5005_ & new_n5604_;
  assign new_n10855_ = new_n5010_ & new_n5610_;
  assign new_n10854_ = new_n5011_ & new_n5611_;
  assign new_n10888_ = new_n5016_ & new_n5617_;
  assign new_n10887_ = new_n5017_ & new_n5618_;
  assign new_n10896_ = new_n5018_ & new_n5619_;
  assign new_n10895_ = new_n5019_ & new_n5620_;
  assign new_n10909_ = new_n5020_ & new_n5622_;
  assign new_n10908_ = new_n5021_ & new_n5623_;
  assign new_n10917_ = new_n5022_ & new_n5624_;
  assign new_n7152_ = ~new_n8696_;
  assign new_n10916_ = new_n5023_ & new_n5625_;
  assign new_n10930_ = new_n5024_ & new_n5627_;
  assign new_n10929_ = new_n5025_ & new_n5628_;
  assign new_n10938_ = new_n5026_ & new_n5629_;
  assign new_n10937_ = new_n5027_ & new_n5630_;
  assign new_n10951_ = new_n5028_ & new_n5632_;
  assign new_n10950_ = new_n5029_ & new_n5633_;
  assign new_n10970_ = new_n5032_ & new_n5636_;
  assign new_n10969_ = new_n5033_ & new_n5637_;
  assign new_n10712_ = new_n11138_ | new_n7424_;
  assign new_n9748_ = new_n10032_ & new_n10033_;
  assign new_n10995_ = new_n5038_ & new_n5642_;
  assign new_n10994_ = new_n5039_ & new_n5643_;
  assign new_n11003_ = new_n5040_ & new_n5644_;
  assign new_n11002_ = new_n5041_ & new_n5645_;
  assign new_n10713_ = new_n7424_ | new_n11137_;
  assign new_n11411_ = new_n5091_ & new_n5700_;
  assign new_n11163_ = new_n7079_ & new_n7061_;
  assign new_n11385_ = new_n5087_ & new_n5696_;
  assign new_n11222_ = new_n7078_ & new_n11231_;
  assign new_n11375_ = new_n5086_ & new_n6632_;
  assign new_n7153_ = ~new_n9748_;
  assign new_n11260_ = new_n7077_ & new_n7060_;
  assign new_n11358_ = new_n5084_ & new_n6630_;
  assign new_n7603_ = new_n7057_ & new_n7252_;
  assign new_n10694_ = new_n4981_ & new_n6620_;
  assign new_n7701_ = new_n5060_ & new_n11151_;
  assign new_n10757_ = new_n10759_ & new_n5588_;
  assign new_n10778_ = new_n10781_ & new_n5593_;
  assign new_n7929_ = new_n4695_ & new_n6481_;
  assign new_n10819_ = new_n10821_ & new_n5602_;
  assign new_n7946_ = new_n4700_ & new_n6484_;
  assign new_n9648_ = new_n10184_ & new_n10185_;
  assign new_n10839_ = new_n10841_ & new_n5607_;
  assign new_n10860_ = new_n10863_ & new_n5612_;
  assign new_n8863_ = new_n7311_ & new_n5301_;
  assign new_n8054_ = new_n6402_ | new_n7440_;
  assign new_n10901_ = new_n10903_ & new_n5621_;
  assign new_n10922_ = new_n10924_ & new_n5626_;
  assign new_n10943_ = new_n10946_ & new_n5631_;
  assign new_n8300_ = new_n5058_ & new_n7701_;
  assign new_n8256_ = new_n4764_ & new_n6536_;
  assign new_n9275_ = new_n9276_ & new_n5370_;
  assign new_n7154_ = ~new_n9648_;
  assign new_n8426_ = new_n4668_ & new_n5226_;
  assign new_n8425_ = new_n4671_ & new_n5228_;
  assign new_n8451_ = new_n4673_ & new_n5230_;
  assign new_n8496_ = new_n4676_ & new_n7560_;
  assign new_n8815_ = new_n4710_ & new_n6493_;
  assign new_n8962_ = new_n4727_ & new_n6508_;
  assign new_n8998_ = new_n7560_ & new_n5324_;
  assign new_n9053_ = new_n4739_ & new_n6518_;
  assign new_n9116_ = new_n4747_ & new_n6524_;
  assign new_n9150_ = new_n7560_ & new_n5349_;
  assign new_n10455_ = new_n7394_ & new_n10586_;
  assign new_n9283_ = new_n4768_ & new_n7039_;
  assign new_n8290_ = new_n7506_ & new_n7155_;
  assign new_n10318_ = new_n4932_ & new_n6610_;
  assign new_n11460_ = new_n5104_ & new_n6639_;
  assign new_n11465_ = new_n5105_ & new_n6640_;
  assign new_n9555_ = new_n4802_ & new_n5390_;
  assign new_n9737_ = new_n9738_ & new_n5419_;
  assign new_n9551_ = new_n4894_ & new_n5493_;
  assign new_n9814_ = new_n9815_ & new_n5431_;
  assign new_n9937_ = new_n9554_ & new_n5453_;
  assign new_n7155_ = ~new_n10455_;
  assign new_n9939_ = new_n4855_ & new_n6593_;
  assign new_n10707_ = new_n4982_ & new_n6621_;
  assign new_n10723_ = new_n4985_ & new_n5581_;
  assign new_n8454_ = new_n6387_ | new_n6425_;
  assign new_n8483_ = new_n6388_ | new_n6426_;
  assign new_n10751_ = new_n4991_ & new_n5587_;
  assign new_n8552_ = new_n6390_ | new_n6428_;
  assign new_n10772_ = new_n4995_ & new_n5592_;
  assign new_n10785_ = new_n4997_ & new_n5595_;
  assign new_n8637_ = new_n6393_ | new_n6431_;
  assign new_n7156_ = ~new_n8867_;
  assign new_n10804_ = new_n5001_ & new_n5599_;
  assign new_n10813_ = new_n5003_ & new_n5601_;
  assign new_n8729_ = new_n6396_ | new_n6434_;
  assign new_n10833_ = new_n5007_ & new_n5606_;
  assign new_n10846_ = new_n5009_ & new_n5609_;
  assign new_n8805_ = new_n6399_ | new_n6437_;
  assign new_n10867_ = new_n5013_ & new_n5614_;
  assign new_n10875_ = new_n5015_ & new_n5616_;
  assign new_n8927_ = new_n6403_ | new_n6441_;
  assign new_n8928_ = new_n6404_ | new_n6442_;
  assign new_n7040_ = ~new_n9120_;
  assign new_n9711_ = new_n10240_ & new_n10241_;
  assign new_n8952_ = new_n6405_ | new_n6443_;
  assign new_n9024_ = new_n6406_ | new_n6444_;
  assign new_n9025_ = new_n6407_ | new_n6445_;
  assign new_n9043_ = new_n6408_ | new_n6446_;
  assign new_n9075_ = new_n6409_ | new_n6447_;
  assign new_n10959_ = new_n5031_ & new_n5635_;
  assign new_n9173_ = new_n6411_ | new_n6449_;
  assign new_n10977_ = new_n5035_ & new_n5639_;
  assign new_n10986_ = new_n5037_ & new_n5641_;
  assign new_n9216_ = new_n6413_ | new_n6451_;
  assign new_n7157_ = ~new_n9711_;
  assign new_n10442_ = new_n6414_ | new_n6452_;
  assign new_n11132_ = new_n5056_ & new_n5660_;
  assign new_n7580_ = new_n11017_ & new_n7390_;
  assign new_n11016_ = IR_REG_0_ & new_n6995_;
  assign new_n11421_ = new_n5093_ & new_n5703_;
  assign new_n7589_ = new_n11017_ & new_n7444_;
  assign new_n11401_ = new_n5090_ & new_n6634_;
  assign new_n11095_ = new_n6207_ & new_n5653_;
  assign new_n11060_ = n1341 & new_n5654_;
  assign new_n11189_ = new_n6213_ & new_n5666_;
  assign new_n9911_ = new_n9945_ & new_n7400_;
  assign new_n11304_ = new_n5070_ & new_n6629_;
  assign new_n11303_ = new_n6223_ & new_n5679_;
  assign new_n10663_ = new_n4970_ & new_n6618_;
  assign new_n7645_ = new_n6007_ & new_n5115_;
  assign new_n10685_ = new_n4978_ & new_n6619_;
  assign new_n7690_ = new_n6010_ & new_n5120_;
  assign new_n11434_ = new_n5100_ & new_n6635_;
  assign new_n7782_ = new_n8416_ & new_n5224_;
  assign new_n7803_ = new_n4580_ & new_n5140_;
  assign new_n7823_ = new_n4583_ & new_n5143_;
  assign new_n7158_ = ~new_n9911_;
  assign new_n7840_ = new_n4586_ & new_n5146_;
  assign new_n7857_ = new_n4589_ & new_n5149_;
  assign new_n7874_ = new_n4592_ & new_n5152_;
  assign new_n7891_ = new_n4595_ & new_n5155_;
  assign new_n7908_ = new_n4598_ & new_n5158_;
  assign new_n7925_ = new_n4601_ & new_n5161_;
  assign new_n7942_ = new_n4604_ & new_n5164_;
  assign new_n7959_ = new_n4607_ & new_n5167_;
  assign new_n7976_ = new_n4610_ & new_n5170_;
  assign new_n7993_ = new_n4613_ & new_n5173_;
  assign new_n7159_ = ~new_n10123_;
  assign new_n8015_ = new_n4969_ & new_n10662_;
  assign new_n8010_ = new_n4616_ & new_n5176_;
  assign new_n8032_ = new_n4967_ & new_n10657_;
  assign new_n8027_ = new_n4619_ & new_n5179_;
  assign new_n8044_ = new_n4622_ & new_n5182_;
  assign new_n8066_ = new_n4972_ & new_n10672_;
  assign new_n8061_ = new_n4625_ & new_n5185_;
  assign new_n8078_ = new_n4628_ & new_n5188_;
  assign new_n8095_ = new_n4631_ & new_n5191_;
  assign new_n8112_ = new_n4634_ & new_n8114_;
  assign new_n8726_ = new_n7243_ & new_n7438_;
  assign new_n8136_ = new_n4959_ & new_n10616_;
  assign new_n8131_ = new_n4637_ & new_n5196_;
  assign new_n8148_ = new_n4640_ & new_n8150_;
  assign new_n8166_ = new_n4643_ & new_n5201_;
  assign new_n8189_ = new_n4960_ & new_n10619_;
  assign new_n8183_ = new_n4646_ & new_n8185_;
  assign new_n8201_ = new_n4649_ & new_n5206_;
  assign new_n7793_ = new_n7418_ | new_n7568_;
  assign new_n8234_ = new_n4655_ & new_n5211_;
  assign new_n8251_ = new_n4658_ & new_n8253_;
  assign new_n7160_ = ~new_n8726_;
  assign new_n8269_ = new_n4661_ & new_n5216_;
  assign new_n8297_ = new_n9235_ & new_n5221_;
  assign new_n7790_ = new_n6379_ | new_n6416_;
  assign new_n8422_ = new_n4672_ & new_n5229_;
  assign new_n8462_ = new_n4674_ & new_n6462_;
  assign new_n8459_ = new_n8474_ & new_n5234_;
  assign new_n8474_ = new_n4675_ & new_n6463_;
  assign new_n8488_ = new_n8504_ & new_n5240_;
  assign new_n8504_ = new_n4678_ & new_n6464_;
  assign new_n8527_ = new_n4681_ & new_n6466_;
  assign new_n7161_ = ~new_n9712_;
  assign new_n8524_ = new_n8537_ & new_n5245_;
  assign new_n8537_ = new_n4682_ & new_n6467_;
  assign new_n8559_ = new_n4683_ & new_n6470_;
  assign new_n8556_ = new_n8565_ & new_n5250_;
  assign new_n8565_ = new_n4684_ & new_n6471_;
  assign new_n8578_ = new_n4685_ & new_n6472_;
  assign new_n8575_ = new_n8587_ & new_n5254_;
  assign new_n8587_ = new_n4686_ & new_n6473_;
  assign new_n8604_ = new_n4688_ & new_n6474_;
  assign new_n8601_ = new_n8630_ & new_n5263_;
  assign new_n9320_ = IR_REG_29_ & new_n7297_;
  assign new_n8630_ = new_n4689_ & new_n6475_;
  assign new_n8645_ = new_n4690_ & new_n6476_;
  assign new_n8642_ = new_n8653_ & new_n5268_;
  assign new_n8653_ = new_n4691_ & new_n6477_;
  assign new_n8680_ = new_n4693_ & new_n6479_;
  assign new_n8677_ = new_n8686_ & new_n5273_;
  assign new_n8686_ = new_n4694_ & new_n6480_;
  assign new_n8704_ = new_n4697_ & new_n6482_;
  assign new_n8701_ = new_n8715_ & new_n5277_;
  assign new_n8715_ = new_n4699_ & new_n6483_;
  assign new_n7162_ = ~new_n9320_;
  assign new_n8737_ = new_n4701_ & new_n6485_;
  assign new_n8734_ = new_n8743_ & new_n5281_;
  assign new_n8743_ = new_n4702_ & new_n6486_;
  assign new_n8756_ = new_n4703_ & new_n6487_;
  assign new_n8753_ = new_n8763_ & new_n5285_;
  assign new_n8763_ = new_n4705_ & new_n6488_;
  assign new_n8783_ = new_n4706_ & new_n6489_;
  assign new_n8780_ = new_n8790_ & new_n5290_;
  assign new_n8790_ = new_n4707_ & new_n6490_;
  assign new_n8811_ = new_n4711_ & new_n6492_;
  assign new_n9057_ = new_n7387_ & new_n7417_;
  assign new_n9470_ = IR_REG_9_ & new_n7287_;
  assign new_n8808_ = new_n8826_ & new_n5295_;
  assign new_n8826_ = new_n4713_ & new_n6494_;
  assign new_n8848_ = new_n4715_ & new_n6496_;
  assign new_n8845_ = new_n8858_ & new_n5300_;
  assign new_n8858_ = new_n4716_ & new_n6497_;
  assign new_n8875_ = new_n4717_ & new_n6498_;
  assign new_n8872_ = new_n8881_ & new_n5305_;
  assign new_n8881_ = new_n4719_ & new_n6499_;
  assign new_n8905_ = new_n4720_ & new_n6501_;
  assign new_n8902_ = new_n8912_ & new_n5310_;
  assign new_n7163_ = ~new_n9470_;
  assign new_n8912_ = new_n4721_ & new_n6502_;
  assign new_n8934_ = new_n4724_ & new_n6505_;
  assign new_n8931_ = new_n8943_ & new_n5314_;
  assign new_n8943_ = new_n4726_ & new_n6506_;
  assign new_n8958_ = new_n4728_ & new_n6507_;
  assign new_n8955_ = new_n8973_ & new_n5320_;
  assign new_n8973_ = new_n4729_ & new_n6509_;
  assign new_n8995_ = new_n4731_ & new_n6511_;
  assign new_n8992_ = new_n9007_ & new_n5326_;
  assign new_n9007_ = new_n4733_ & new_n6512_;
  assign new_n9382_ = IR_REG_21_ & new_n7296_;
  assign new_n9031_ = new_n4736_ & new_n6515_;
  assign new_n9028_ = new_n9037_ & new_n5331_;
  assign new_n9037_ = new_n4737_ & new_n6516_;
  assign new_n9049_ = new_n4740_ & new_n6517_;
  assign new_n9046_ = new_n9064_ & new_n5335_;
  assign new_n9064_ = new_n4742_ & new_n6519_;
  assign new_n9084_ = new_n4743_ & new_n6520_;
  assign new_n9081_ = new_n9092_ & new_n5340_;
  assign new_n9092_ = new_n4744_ & new_n6521_;
  assign new_n9112_ = new_n4748_ & new_n6523_;
  assign new_n7164_ = ~new_n9382_;
  assign new_n9109_ = new_n9127_ & new_n5345_;
  assign new_n9127_ = new_n4750_ & new_n6525_;
  assign new_n9147_ = new_n4752_ & new_n6527_;
  assign new_n9144_ = new_n9157_ & new_n5350_;
  assign new_n9157_ = new_n4753_ & new_n6528_;
  assign new_n9179_ = new_n4756_ & new_n6530_;
  assign new_n9176_ = new_n9186_ & new_n5354_;
  assign new_n9186_ = new_n4757_ & new_n6531_;
  assign new_n9202_ = new_n4759_ & new_n6532_;
  assign new_n9199_ = new_n9209_ & new_n5358_;
  assign new_n9367_ = IR_REG_23_ & new_n7283_;
  assign new_n9209_ = new_n4760_ & new_n6533_;
  assign new_n9222_ = new_n4762_ & new_n6534_;
  assign new_n9219_ = new_n9229_ & new_n5362_;
  assign new_n9229_ = new_n4763_ & new_n6535_;
  assign new_n9250_ = new_n4765_ & new_n6537_;
  assign new_n9247_ = new_n9257_ & new_n5366_;
  assign new_n9257_ = new_n4766_ & new_n6538_;
  assign new_n8398_ = new_n6381_ | new_n6421_;
  assign new_n9267_ = new_n9235_ & new_n5368_;
  assign new_n9336_ = new_n7313_ | IR_REG_26_;
  assign new_n7165_ = ~new_n9367_;
  assign new_n9389_ = new_n7308_ | IR_REG_19_;
  assign new_n9403_ = new_n7309_ | IR_REG_17_;
  assign new_n9485_ = IR_REG_7_ & new_n7001_;
  assign new_n9506_ = new_n7404_ | IR_REG_3_;
  assign new_n9523_ = IR_REG_2_ & new_n7002_;
  assign new_n9543_ = new_n4801_ & new_n5388_;
  assign new_n9541_ = new_n9549_ & new_n5389_;
  assign new_n9571_ = new_n4803_ & new_n5392_;
  assign new_n9569_ = new_n9575_ & new_n5393_;
  assign new_n9575_ = new_n4804_ & new_n6570_;
  assign new_n8669_ = new_n7241_ & new_n7509_;
  assign new_n9586_ = new_n4805_ & new_n5394_;
  assign new_n9584_ = new_n9589_ & new_n5395_;
  assign new_n9589_ = new_n4806_ & new_n6571_;
  assign new_n9600_ = new_n4807_ & new_n5397_;
  assign new_n9598_ = new_n9604_ & new_n5398_;
  assign new_n9604_ = new_n4808_ & new_n6572_;
  assign new_n9615_ = new_n4809_ & new_n5399_;
  assign new_n9613_ = new_n9619_ & new_n5400_;
  assign new_n9619_ = new_n4810_ & new_n6573_;
  assign new_n9627_ = new_n9633_ & new_n5402_;
  assign new_n7166_ = ~new_n8669_;
  assign new_n9633_ = new_n4812_ & new_n6574_;
  assign new_n9651_ = new_n4813_ & new_n5403_;
  assign new_n9649_ = new_n9654_ & new_n5404_;
  assign new_n9654_ = new_n4814_ & new_n6576_;
  assign new_n9665_ = new_n4815_ & new_n5406_;
  assign new_n9663_ = new_n9669_ & new_n5407_;
  assign new_n9669_ = new_n4822_ & new_n6577_;
  assign new_n9700_ = new_n4823_ & new_n5412_;
  assign new_n9698_ = new_n9704_ & new_n5413_;
  assign new_n9704_ = new_n4824_ & new_n6579_;
  assign new_n8697_ = new_n7242_ & new_n7385_;
  assign new_n9713_ = new_n9717_ & new_n5415_;
  assign new_n9717_ = new_n4826_ & new_n6580_;
  assign new_n9729_ = new_n4827_ & new_n5417_;
  assign new_n9727_ = new_n9733_ & new_n5418_;
  assign new_n9751_ = new_n4829_ & new_n5420_;
  assign new_n9749_ = new_n9755_ & new_n5421_;
  assign new_n9755_ = new_n4830_ & new_n6581_;
  assign new_n9765_ = new_n4831_ & new_n5423_;
  assign new_n9763_ = new_n9769_ & new_n5424_;
  assign new_n9769_ = new_n4832_ & new_n6582_;
  assign new_n7167_ = ~new_n8697_;
  assign new_n9780_ = new_n4833_ & new_n5425_;
  assign new_n9778_ = new_n9783_ & new_n5426_;
  assign new_n9783_ = new_n4834_ & new_n6583_;
  assign new_n9793_ = new_n4835_ & new_n5427_;
  assign new_n9791_ = new_n9797_ & new_n5428_;
  assign new_n9797_ = new_n4836_ & new_n6584_;
  assign new_n9807_ = new_n4837_ & new_n5429_;
  assign new_n9805_ = new_n9810_ & new_n5430_;
  assign new_n9826_ = new_n4839_ & new_n5433_;
  assign new_n9824_ = new_n9830_ & new_n5434_;
  assign new_n7041_ = ~new_n9057_;
  assign new_n7168_ = ~new_n9242_;
  assign new_n9830_ = new_n4840_ & new_n6585_;
  assign new_n9841_ = new_n4841_ & new_n5435_;
  assign new_n9839_ = new_n9845_ & new_n5436_;
  assign new_n9845_ = new_n4842_ & new_n6586_;
  assign new_n9856_ = new_n4843_ & new_n5437_;
  assign new_n9854_ = new_n9860_ & new_n5438_;
  assign new_n9860_ = new_n4844_ & new_n6587_;
  assign new_n9869_ = new_n4846_ & new_n5440_;
  assign new_n9878_ = new_n4847_ & new_n5442_;
  assign new_n9876_ = new_n9882_ & new_n5443_;
  assign new_n10159_ = new_n9681_ & new_n8083_;
  assign new_n9882_ = new_n4848_ & new_n6588_;
  assign new_n9890_ = new_n4849_ & new_n5444_;
  assign new_n9888_ = new_n9893_ & new_n5445_;
  assign new_n9893_ = new_n4851_ & new_n6589_;
  assign new_n9915_ = new_n4852_ & new_n5449_;
  assign new_n9913_ = new_n9919_ & new_n5450_;
  assign new_n9919_ = new_n4853_ & new_n6591_;
  assign new_n9930_ = new_n4854_ & new_n5451_;
  assign new_n9928_ = new_n9934_ & new_n5452_;
  assign new_n9934_ = new_n4856_ & new_n6592_;
  assign new_n7169_ = ~new_n10159_;
  assign new_n9949_ = new_n9953_ & new_n5456_;
  assign new_n9953_ = new_n4858_ & new_n6594_;
  assign new_n9961_ = new_n4859_ & new_n5457_;
  assign new_n9959_ = new_n9964_ & new_n5458_;
  assign new_n9964_ = new_n4860_ & new_n6595_;
  assign new_n9975_ = new_n4861_ & new_n5459_;
  assign new_n9973_ = new_n9979_ & new_n5460_;
  assign new_n9979_ = new_n4862_ & new_n6596_;
  assign new_n9989_ = new_n4863_ & new_n5463_;
  assign new_n9987_ = new_n9993_ & new_n5464_;
  assign new_n9425_ = IR_REG_15_ & new_n7284_;
  assign new_n9993_ = new_n4892_ & new_n6597_;
  assign new_n10104_ = new_n4893_ & new_n5491_;
  assign new_n10102_ = new_n10110_ & new_n5492_;
  assign new_n10110_ = new_n4929_ & new_n6604_;
  assign new_n10329_ = new_n4937_ & new_n6611_;
  assign new_n8419_ = new_n10707_ & new_n5578_;
  assign new_n8429_ = new_n10717_ & new_n5579_;
  assign new_n10717_ = new_n4983_ & new_n6622_;
  assign new_n10724_ = new_n4984_ & new_n5580_;
  assign new_n10752_ = new_n4990_ & new_n5586_;
  assign new_n7170_ = ~new_n9425_;
  assign new_n10773_ = new_n4994_ & new_n5591_;
  assign new_n10786_ = new_n4996_ & new_n5594_;
  assign new_n10805_ = new_n5000_ & new_n5598_;
  assign new_n10814_ = new_n5002_ & new_n5600_;
  assign new_n10834_ = new_n5006_ & new_n5605_;
  assign new_n10847_ = new_n5008_ & new_n5608_;
  assign new_n10868_ = new_n5012_ & new_n5613_;
  assign new_n10876_ = new_n5014_ & new_n5615_;
  assign new_n10960_ = new_n5030_ & new_n5634_;
  assign new_n10978_ = new_n5034_ & new_n5638_;
  assign new_n9440_ = IR_REG_13_ & new_n7285_;
  assign new_n10987_ = new_n5036_ & new_n5640_;
  assign new_n11133_ = new_n5055_ & new_n5659_;
  assign new_n11011_ = new_n5042_ & new_n5646_;
  assign new_n11028_ = new_n5044_ & new_n6623_;
  assign new_n11025_ = new_n5043_ & new_n5647_;
  assign new_n11042_ = new_n5045_ & new_n5649_;
  assign new_n11040_ = new_n5046_ & new_n7112_;
  assign new_n11061_ = new_n5047_ & new_n5651_;
  assign new_n11083_ = new_n5048_ & new_n5652_;
  assign new_n11081_ = new_n5061_ & new_n7112_;
  assign new_n7171_ = ~new_n9440_;
  assign new_n11154_ = new_n5062_ & new_n5663_;
  assign new_n11174_ = new_n5063_ & new_n5665_;
  assign new_n11195_ = new_n5064_ & new_n5668_;
  assign new_n11214_ = new_n5065_ & new_n5670_;
  assign new_n11233_ = new_n5066_ & new_n5672_;
  assign new_n11252_ = new_n5067_ & new_n5674_;
  assign new_n11271_ = new_n5068_ & new_n5676_;
  assign new_n11291_ = new_n5069_ & new_n5678_;
  assign new_n7570_ = new_n4556_ & new_n5108_;
  assign new_n7592_ = new_n4557_ & new_n5110_;
  assign new_n9455_ = IR_REG_11_ & new_n7286_;
  assign new_n7611_ = new_n4558_ & new_n5112_;
  assign new_n7630_ = new_n4559_ & new_n5114_;
  assign new_n7651_ = new_n4560_ & new_n5117_;
  assign new_n7673_ = new_n4561_ & new_n5119_;
  assign new_n7695_ = new_n4562_ & new_n5122_;
  assign new_n7768_ = new_n4576_ & new_n7104_;
  assign new_n7776_ = new_n4578_ & new_n7104_;
  assign new_n7784_ = new_n7791_ & new_n5139_;
  assign new_n7791_ = new_n4579_ & new_n6459_;
  assign new_n7810_ = new_n4582_ & new_n5142_;
  assign new_n7172_ = ~new_n9455_;
  assign new_n7811_ = new_n4581_ & new_n5141_;
  assign new_n7829_ = new_n4585_ & new_n5145_;
  assign new_n7830_ = new_n4584_ & new_n5144_;
  assign new_n7846_ = new_n4588_ & new_n5148_;
  assign new_n7847_ = new_n4587_ & new_n5147_;
  assign new_n7863_ = new_n4591_ & new_n5151_;
  assign new_n7864_ = new_n4590_ & new_n5150_;
  assign new_n7880_ = new_n4594_ & new_n5154_;
  assign new_n7881_ = new_n4593_ & new_n5153_;
  assign new_n7897_ = new_n4597_ & new_n5157_;
  assign new_n7173_ = ~new_n9523_;
  assign new_n7898_ = new_n4596_ & new_n5156_;
  assign new_n7914_ = new_n4600_ & new_n5160_;
  assign new_n7915_ = new_n4599_ & new_n5159_;
  assign new_n7931_ = new_n4603_ & new_n5163_;
  assign new_n7932_ = new_n4602_ & new_n5162_;
  assign new_n7948_ = new_n4606_ & new_n5166_;
  assign new_n7949_ = new_n4605_ & new_n5165_;
  assign new_n7965_ = new_n4609_ & new_n5169_;
  assign new_n7966_ = new_n4608_ & new_n5168_;
  assign new_n7982_ = new_n4612_ & new_n5172_;
  assign new_n8824_ = new_n7452_ & new_n7478_;
  assign new_n7174_ = ~new_n9485_;
  assign new_n7983_ = new_n4611_ & new_n5171_;
  assign new_n7999_ = new_n4615_ & new_n5175_;
  assign new_n8000_ = new_n4614_ & new_n5174_;
  assign new_n8016_ = new_n4618_ & new_n5178_;
  assign new_n8017_ = new_n4617_ & new_n5177_;
  assign new_n8033_ = new_n4621_ & new_n5181_;
  assign new_n8034_ = new_n4620_ & new_n5180_;
  assign new_n8050_ = new_n4624_ & new_n5184_;
  assign new_n8051_ = new_n4623_ & new_n5183_;
  assign new_n8067_ = new_n4627_ & new_n5187_;
  assign new_n7175_ = ~new_n10174_;
  assign new_n8068_ = new_n4626_ & new_n5186_;
  assign new_n8084_ = new_n4630_ & new_n5190_;
  assign new_n8085_ = new_n4629_ & new_n5189_;
  assign new_n8101_ = new_n4633_ & new_n5193_;
  assign new_n8102_ = new_n4632_ & new_n5192_;
  assign new_n8120_ = new_n4636_ & new_n5195_;
  assign new_n8121_ = new_n4635_ & new_n5194_;
  assign new_n8137_ = new_n4639_ & new_n5198_;
  assign new_n8138_ = new_n4638_ & new_n5197_;
  assign new_n8155_ = new_n4642_ & new_n5200_;
  assign new_n7176_ = ~new_n7782_;
  assign new_n8156_ = new_n4641_ & new_n5199_;
  assign new_n8172_ = new_n4645_ & new_n5203_;
  assign new_n8173_ = new_n4644_ & new_n5202_;
  assign new_n8190_ = new_n4648_ & new_n5205_;
  assign new_n8191_ = new_n4647_ & new_n5204_;
  assign new_n8207_ = new_n4651_ & new_n5208_;
  assign new_n8208_ = new_n4650_ & new_n5207_;
  assign new_n8224_ = new_n4654_ & new_n5210_;
  assign new_n8225_ = new_n4653_ & new_n5209_;
  assign new_n8218_ = new_n4652_ & new_n8220_;
  assign new_n8518_ = new_n7845_ & new_n8553_;
  assign new_n8240_ = new_n4657_ & new_n5213_;
  assign new_n8241_ = new_n4656_ & new_n5212_;
  assign new_n8258_ = new_n4660_ & new_n5215_;
  assign new_n8259_ = new_n4659_ & new_n5214_;
  assign new_n8275_ = new_n4663_ & new_n5218_;
  assign new_n8276_ = new_n4662_ & new_n5217_;
  assign new_n8282_ = new_n8293_ & new_n5220_;
  assign new_n8293_ = new_n4665_ & new_n6461_;
  assign new_n8303_ = new_n8402_ & new_n5222_;
  assign new_n8307_ = new_n4666_ & new_n5223_;
  assign new_n7177_ = ~new_n8518_;
  assign new_n8423_ = new_n7200_ & new_n5225_;
  assign new_n8460_ = new_n7819_ & new_n5231_;
  assign new_n8489_ = new_n7836_ & new_n5237_;
  assign new_n8525_ = new_n7853_ & new_n5242_;
  assign new_n8557_ = new_n7870_ & new_n5248_;
  assign new_n8576_ = new_n7887_ & new_n5252_;
  assign new_n8602_ = new_n7904_ & new_n5257_;
  assign new_n8643_ = new_n7921_ & new_n5265_;
  assign new_n8678_ = new_n7938_ & new_n5271_;
  assign new_n8702_ = new_n7955_ & new_n5274_;
  assign new_n8513_ = new_n7391_ & new_n7454_;
  assign new_n8735_ = new_n7972_ & new_n5279_;
  assign new_n8754_ = new_n7989_ & new_n5283_;
  assign new_n8781_ = new_n8006_ & new_n5288_;
  assign new_n8809_ = new_n8023_ & new_n5292_;
  assign new_n8846_ = new_n8040_ & new_n5297_;
  assign new_n8873_ = new_n8057_ & new_n5303_;
  assign new_n8903_ = new_n8074_ & new_n5308_;
  assign new_n8932_ = new_n8091_ & new_n5312_;
  assign new_n8956_ = new_n8108_ & new_n5317_;
  assign new_n8993_ = new_n8127_ & new_n5322_;
  assign new_n7178_ = ~new_n8513_;
  assign new_n9029_ = new_n8144_ & new_n5329_;
  assign new_n9047_ = new_n8162_ & new_n5333_;
  assign new_n9082_ = new_n8179_ & new_n5338_;
  assign new_n9110_ = new_n8197_ & new_n5343_;
  assign new_n9145_ = new_n8214_ & new_n5347_;
  assign new_n9177_ = new_n8230_ & new_n5352_;
  assign new_n9200_ = new_n8247_ & new_n5356_;
  assign new_n9220_ = new_n8265_ & new_n5360_;
  assign new_n9248_ = new_n8281_ & new_n5364_;
  assign new_n8397_ = new_n9263_ & new_n5367_;
  assign new_n8666_ = new_n7244_ & new_n7456_;
  assign new_n9263_ = new_n4767_ & new_n6539_;
  assign new_n9309_ = IR_REG_30_ & new_n5371_;
  assign new_n9325_ = IR_REG_28_ & new_n5372_;
  assign new_n9333_ = IR_REG_27_ & new_n5373_;
  assign new_n9347_ = IR_REG_25_ & new_n5374_;
  assign new_n9356_ = IR_REG_24_ & new_n5375_;
  assign new_n9371_ = IR_REG_22_ & new_n5376_;
  assign new_n9386_ = IR_REG_20_ & new_n5377_;
  assign new_n9395_ = new_n4780_ & new_n9313_;
  assign new_n9400_ = IR_REG_18_ & new_n5378_;
  assign new_n7179_ = ~new_n8666_;
  assign new_n9409_ = new_n4783_ & new_n9313_;
  assign new_n9414_ = IR_REG_16_ & new_n5379_;
  assign new_n9429_ = IR_REG_14_ & new_n5380_;
  assign new_n9444_ = IR_REG_12_ & new_n5381_;
  assign new_n9459_ = IR_REG_10_ & new_n5382_;
  assign new_n9474_ = IR_REG_8_ & new_n5383_;
  assign new_n9489_ = IR_REG_6_ & new_n5384_;
  assign new_n9503_ = IR_REG_4_ & new_n5385_;
  assign new_n9512_ = IR_REG_3_ & new_n5386_;
  assign new_n9527_ = IR_REG_1_ & new_n5387_;
  assign new_n8896_ = new_n8066_ & new_n8927_;
  assign new_n9570_ = new_n9571_ & new_n5391_;
  assign new_n9599_ = new_n9600_ & new_n5396_;
  assign new_n9628_ = new_n9629_ & new_n5401_;
  assign new_n9664_ = new_n9665_ & new_n5405_;
  assign new_n9714_ = new_n4825_ & new_n5414_;
  assign new_n9728_ = new_n9729_ & new_n5416_;
  assign new_n9764_ = new_n9765_ & new_n5422_;
  assign new_n9825_ = new_n9826_ & new_n5432_;
  assign new_n9870_ = new_n4845_ & new_n5439_;
  assign new_n9877_ = new_n9878_ & new_n5441_;
  assign new_n7042_ = ~new_n8824_;
  assign new_n7180_ = ~new_n8896_;
  assign new_n9914_ = new_n9915_ & new_n5448_;
  assign new_n9950_ = new_n4857_ & new_n5455_;
  assign new_n9988_ = new_n9989_ & new_n5462_;
  assign new_n11041_ = new_n11042_ & new_n5648_;
  assign new_n11062_ = new_n7199_ & new_n5650_;
  assign new_n11155_ = new_n7136_ & new_n5662_;
  assign new_n11175_ = new_n7137_ & new_n5664_;
  assign new_n11196_ = new_n7138_ & new_n5667_;
  assign new_n11215_ = new_n7139_ & new_n5669_;
  assign new_n11234_ = new_n7140_ & new_n5671_;
  assign new_n7181_ = ~new_n8116_;
  assign new_n11253_ = new_n7141_ & new_n5673_;
  assign new_n11272_ = new_n7142_ & new_n5675_;
  assign new_n11292_ = new_n7143_ & new_n5677_;
  assign new_n7571_ = new_n7131_ & new_n5107_;
  assign new_n7593_ = new_n7127_ & new_n5109_;
  assign new_n7612_ = new_n7133_ & new_n5111_;
  assign new_n7631_ = new_n7129_ & new_n5113_;
  assign new_n7652_ = new_n7130_ & new_n5116_;
  assign new_n7674_ = new_n7132_ & new_n5118_;
  assign new_n7696_ = new_n7128_ & new_n5121_;
  assign new_n8986_ = new_n8119_ & new_n9024_;
  assign new_n7769_ = new_n4575_ & new_n5136_;
  assign new_n7777_ = new_n4577_ & new_n5137_;
  assign new_n7785_ = new_n7786_ & new_n5138_;
  assign new_n8283_ = new_n8284_ & new_n5219_;
  assign new_n9306_ = new_n4769_ & new_n6540_;
  assign new_n9315_ = new_n4770_ & new_n6541_;
  assign new_n9322_ = new_n4771_ & new_n6542_;
  assign new_n9330_ = new_n4772_ & new_n6543_;
  assign new_n9339_ = new_n4773_ & new_n6544_;
  assign new_n9344_ = new_n4774_ & new_n6545_;
  assign new_n7182_ = ~new_n8986_;
  assign new_n9353_ = new_n4775_ & new_n6546_;
  assign new_n9362_ = new_n4776_ & new_n6547_;
  assign new_n9368_ = new_n4777_ & new_n6548_;
  assign new_n9377_ = new_n4778_ & new_n6549_;
  assign new_n9383_ = new_n4779_ & new_n6550_;
  assign new_n9392_ = new_n4781_ & new_n6551_;
  assign new_n9397_ = new_n4782_ & new_n6552_;
  assign new_n9406_ = new_n4784_ & new_n6553_;
  assign new_n9411_ = new_n4785_ & new_n6554_;
  assign new_n9420_ = new_n4786_ & new_n6555_;
  assign new_n7183_ = ~new_n8151_;
  assign new_n9426_ = new_n4787_ & new_n6556_;
  assign new_n9435_ = new_n4788_ & new_n6557_;
  assign new_n9441_ = new_n4789_ & new_n6558_;
  assign new_n9450_ = new_n4790_ & new_n6559_;
  assign new_n9456_ = new_n4791_ & new_n6560_;
  assign new_n9465_ = new_n4792_ & new_n6561_;
  assign new_n9471_ = new_n4793_ & new_n6562_;
  assign new_n9479_ = new_n4794_ & new_n6563_;
  assign new_n9486_ = new_n4795_ & new_n6564_;
  assign new_n9495_ = new_n4796_ & new_n6565_;
  assign new_n7184_ = ~new_n8186_;
  assign new_n9500_ = new_n4797_ & new_n6566_;
  assign new_n9509_ = new_n4798_ & new_n6567_;
  assign new_n9517_ = new_n4799_ & new_n6568_;
  assign new_n9524_ = new_n4800_ & new_n6569_;
  assign new_n8750_ = new_n6397_ | new_n6435_;
  assign new_n8100_ = new_n4966_ & new_n10651_;
  assign new_n8774_ = new_n6398_ | new_n6436_;
  assign new_n8521_ = new_n6391_ | new_n6429_;
  assign new_n8869_ = new_n6401_ | new_n6439_;
  assign new_n8553_ = new_n6389_ | new_n6427_;
  assign new_n8221_ = new_n9172_ & new_n9192_;
  assign new_n8674_ = new_n6394_ | new_n6432_;
  assign new_n8841_ = new_n6400_ | new_n6438_;
  assign new_n9106_ = new_n6410_ | new_n6448_;
  assign new_n9171_ = new_n6412_ | new_n6450_;
  assign new_n8728_ = new_n6395_ | new_n6433_;
  assign new_n8206_ = new_n4956_ & new_n10608_;
  assign new_n7964_ = new_n4979_ & new_n10691_;
  assign new_n8596_ = new_n6392_ | new_n6430_;
  assign new_n8257_ = new_n4954_ & new_n10595_;
  assign new_n8154_ = new_n4957_ & new_n10610_;
  assign new_n7185_ = ~new_n8221_;
  assign new_n8119_ = new_n4965_ & new_n10648_;
  assign new_n10586_ = new_n6415_ | new_n6453_;
  assign new_n9278_ = new_n11441_ & new_n7283_;
  assign new_n11036_ = new_n11428_ | new_n6456_;
  assign new_n11417_ = new_n5092_ & new_n5702_;
  assign new_n9166_ = new_n4758_ & new_n5355_;
  assign new_n8794_ = new_n4712_ & new_n8862_;
  assign new_n8916_ = new_n4725_ & new_n8117_;
  assign new_n8152_ = new_n4741_ & new_n8187_;
  assign new_n11066_ = new_n7483_ | new_n6455_;
  assign new_n7186_ = ~new_n8254_;
  assign new_n10531_ = new_n4961_ & new_n5562_;
  assign new_n10033_ = new_n4873_ & new_n5474_;
  assign new_n10054_ = new_n4877_ & new_n5477_;
  assign new_n10095_ = new_n4890_ & new_n5489_;
  assign new_n10185_ = new_n4901_ & new_n5502_;
  assign new_n10195_ = new_n4904_ & new_n5506_;
  assign new_n10241_ = new_n4916_ & new_n5517_;
  assign new_n10164_ = new_n4920_ & new_n5521_;
  assign new_n10042_ = new_n4885_ & new_n5485_;
  assign new_n10005_ = new_n4865_ & new_n5465_;
  assign new_n7187_ = ~new_n10121_;
  assign new_n10063_ = new_n4879_ & new_n5480_;
  assign new_n10208_ = new_n4906_ & new_n5508_;
  assign new_n10228_ = new_n4914_ & new_n5515_;
  assign new_n10150_ = new_n4924_ & new_n5525_;
  assign new_n10219_ = new_n4912_ & new_n5513_;
  assign new_n11114_ = new_n7451_ & new_n5657_;
  assign new_n7981_ = new_n4977_ & new_n10684_;
  assign new_n8239_ = new_n4955_ & new_n10598_;
  assign new_n10703_ = new_n5103_ & new_n7450_;
  assign new_n7722_ = new_n7096_ & new_n5126_;
  assign new_n8971_ = new_n7458_ & new_n7281_;
  assign new_n10158_ = new_n11114_ & new_n8928_;
  assign new_n9265_ = new_n11451_ & new_n7297_;
  assign new_n8731_ = new_n7179_ & new_n5282_;
  assign new_n8690_ = new_n4698_ & new_n8747_;
  assign new_n9300_ = new_n10318_ & new_n7260_;
  assign new_n8551_ = new_n7178_ & new_n5251_;
  assign new_n8572_ = new_n4687_ & new_n5256_;
  assign new_n11017_ = new_n5101_ & new_n6999_;
  assign new_n10596_ = new_n5094_ & new_n5704_;
  assign new_n7689_ = new_n10685_ & new_n7308_;
  assign new_n9775_ = new_n4868_ & new_n5467_;
  assign new_n7188_ = ~new_n10158_;
  assign new_n8444_ = new_n6978_ & new_n5233_;
  assign new_n8891_ = new_n4730_ & new_n5321_;
  assign new_n9133_ = new_n7507_ | new_n6419_;
  assign new_n9944_ = new_n4922_ & new_n5523_;
  assign new_n10649_ = new_n11358_ & new_n7286_;
  assign new_n10611_ = new_n11375_ & new_n7287_;
  assign new_n7646_ = new_n10663_ & new_n7309_;
  assign new_n7609_ = REG1_REG_14_ & new_n5128_;
  assign new_n8468_ = new_n7462_ & new_n5547_;
  assign new_n10378_ = new_n7302_ & new_n5570_;
  assign new_n7189_ = ~new_n7581_;
  assign new_n7819_ = new_n8462_ & new_n5232_;
  assign new_n7836_ = new_n8491_ & new_n5238_;
  assign new_n7853_ = new_n8527_ & new_n5243_;
  assign new_n7870_ = new_n8559_ & new_n5249_;
  assign new_n7887_ = new_n8578_ & new_n5253_;
  assign new_n7904_ = new_n8604_ & new_n5258_;
  assign new_n7921_ = new_n8645_ & new_n5266_;
  assign new_n7938_ = new_n8680_ & new_n5272_;
  assign new_n7955_ = new_n8704_ & new_n5275_;
  assign new_n7972_ = new_n8737_ & new_n5280_;
  assign new_n7190_ = ~new_n7603_;
  assign new_n7989_ = new_n8756_ & new_n5284_;
  assign new_n8006_ = new_n8783_ & new_n5289_;
  assign new_n8023_ = new_n8811_ & new_n5293_;
  assign new_n8040_ = new_n8848_ & new_n5298_;
  assign new_n8057_ = new_n8875_ & new_n5304_;
  assign new_n8074_ = new_n8905_ & new_n5309_;
  assign new_n8091_ = new_n8934_ & new_n5313_;
  assign new_n8108_ = new_n8958_ & new_n5318_;
  assign new_n8127_ = new_n8995_ & new_n5323_;
  assign new_n8144_ = new_n9031_ & new_n5330_;
  assign new_n7191_ = ~new_n7621_;
  assign new_n8162_ = new_n9049_ & new_n5334_;
  assign new_n8179_ = new_n9084_ & new_n5339_;
  assign new_n8197_ = new_n9112_ & new_n5344_;
  assign new_n8214_ = new_n9147_ & new_n5348_;
  assign new_n8230_ = new_n9179_ & new_n5353_;
  assign new_n8247_ = new_n9202_ & new_n5357_;
  assign new_n8265_ = new_n9222_ & new_n5361_;
  assign new_n8281_ = new_n9250_ & new_n5365_;
  assign new_n8667_ = new_n8770_ & new_n5287_;
  assign new_n8981_ = new_n9071_ & new_n5337_;
  assign new_n7192_ = ~new_n11070_;
  assign new_n7657_ = new_n4975_ & new_n10679_;
  assign new_n8304_ = new_n8399_ & new_n7059_;
  assign new_n8115_ = new_n4664_ & new_n8413_;
  assign new_n9554_ = new_n10127_ & new_n7230_;
  assign new_n8171_ = new_n4958_ & new_n10613_;
  assign new_n7998_ = new_n4974_ & new_n10677_;
  assign new_n9235_ = new_n11130_ & new_n5658_;
  assign new_n8083_ = new_n4971_ & new_n10670_;
  assign new_n8049_ = new_n4980_ & new_n10693_;
  assign new_n9293_ = new_n10703_ & new_n7410_;
  assign new_n7193_ = ~new_n11163_;
  assign new_n8274_ = new_n4952_ & new_n10589_;
  assign new_n7798_ = new_n7568_ | new_n7196_;
  assign new_n8291_ = new_n9272_ & new_n5369_;
  assign new_n10122_ = new_n7386_ | new_n7215_;
  assign new_n11159_ = new_n5089_ & new_n5698_;
  assign new_n11106_ = new_n11446_ & new_n7000_;
  assign new_n8536_ = new_n10489_ & new_n5549_;
  assign new_n9948_ = new_n10166_ & new_n5500_;
  assign new_n9905_ = new_n9909_ & new_n5447_;
  assign new_n9821_ = new_n10065_ & new_n5479_;
  assign new_n7194_ = ~new_n11222_;
  assign new_n9745_ = new_n10044_ & new_n5476_;
  assign new_n9567_ = new_n9803_ & new_n5461_;
  assign new_n9986_ = new_n10178_ & new_n5501_;
  assign new_n11090_ = new_n11079_ & new_n5699_;
  assign new_n11248_ = new_n11231_ & new_n5693_;
  assign new_n8968_ = new_n8119_ & new_n7249_;
  assign new_n10652_ = new_n5082_ & new_n11351_;
  assign new_n8472_ = new_n7232_ & new_n7828_;
  assign new_n10319_ = new_n5106_ & new_n5706_;
  assign new_n8899_ = new_n4723_ & new_n7058_;
  assign new_n7195_ = ~new_n11260_;
  assign new_n9432_ = new_n7285_ | IR_REG_13_;
  assign new_n9447_ = new_n7286_ | IR_REG_11_;
  assign new_n9417_ = new_n7284_ | IR_REG_15_;
  assign new_n10119_ = new_n5102_ & new_n11457_;
  assign new_n10138_ = new_n5053_ & new_n11129_;
  assign new_n8969_ = new_n7475_ & new_n5325_;
  assign new_n8629_ = new_n8674_ & new_n7509_;
  assign new_n8854_ = new_n7382_ & new_n8869_;
  assign new_n10411_ = new_n7235_ & new_n8015_;
  assign new_n9646_ = new_n7075_ & new_n5504_;
  assign new_n10279_ = new_n8450_ & new_n7550_;
  assign new_n10415_ = new_n7981_ & new_n7244_;
  assign new_n9492_ = new_n7276_ | IR_REG_5_;
  assign new_n10375_ = new_n8100_ & new_n7248_;
  assign new_n8615_ = new_n8637_ & new_n7395_;
  assign new_n8512_ = new_n7070_ & new_n7094_;
  assign new_n7617_ = new_n4968_ & new_n10659_;
  assign new_n7576_ = new_n4973_ & new_n10674_;
  assign new_n7605_ = new_n10694_ & new_n7284_;
  assign new_n10614_ = new_n5095_ & new_n5705_;
  assign new_n10617_ = new_n5085_ & new_n11366_;
  assign new_n7043_ = ~new_n8971_;
  assign new_n7196_ = ~new_n10279_;
  assign new_n10464_ = new_n8083_ & new_n7247_;
  assign new_n8413_ = new_n7118_ & new_n7550_;
  assign new_n7772_ = new_n10703_ & new_n5532_;
  assign new_n8747_ = new_n4704_ & new_n8794_;
  assign new_n8862_ = new_n4718_ & new_n8916_;
  assign new_n8117_ = new_n4732_ & new_n8152_;
  assign new_n8187_ = new_n4749_ & new_n7429_;
  assign new_n11179_ = new_n11432_ | new_n6454_;
  assign new_n8822_ = new_n7515_ & new_n5299_;
  assign new_n7738_ = new_n11347_ & new_n5691_;
  assign new_n7197_ = ~new_n9091_;
  assign new_n10416_ = new_n7947_ & new_n7242_;
  assign new_n8989_ = new_n4735_ & new_n7125_;
  assign new_n8502_ = new_n8553_ & new_n7447_;
  assign new_n9126_ = new_n7525_ & new_n7151_;
  assign new_n8614_ = new_n7482_ & new_n7259_;
  assign new_n8399_ = new_n7076_ & new_n10317_;
  assign new_n9282_ = new_n5096_ & new_n11439_;
  assign new_n10635_ = new_n7444_ & new_n7390_;
  assign new_n9685_ = new_n11116_ & new_n7066_;
  assign new_n8407_ = new_n7059_ & new_n7386_;
  assign new_n7198_ = ~new_n8941_;
  assign new_n9122_ = new_n7237_ & new_n8206_;
  assign new_n9059_ = new_n7371_ & new_n8171_;
  assign new_n9359_ = new_n7283_ | IR_REG_23_;
  assign new_n9374_ = new_n7296_ | IR_REG_21_;
  assign new_n9462_ = new_n7287_ | IR_REG_9_;
  assign new_n7739_ = new_n11304_ & new_n7285_;
  assign new_n10593_ = new_n7276_ & new_n11401_;
  assign new_n7574_ = new_n7576_ & new_n5708_;
  assign new_n4556_ = ~new_n7574_;
  assign new_n7596_ = new_n6003_ & new_n7455_;
  assign new_n9632_ = REG3_REG_3_ & n1332;
  assign new_n4557_ = ~new_n7596_;
  assign new_n7615_ = new_n7617_ & new_n5711_;
  assign new_n4558_ = ~new_n7615_;
  assign new_n7634_ = new_n6006_ & new_n7513_;
  assign new_n4559_ = ~new_n7634_;
  assign new_n7655_ = new_n7657_ & new_n5716_;
  assign new_n4560_ = ~new_n7655_;
  assign new_n7677_ = new_n6009_ & new_n7537_;
  assign new_n4561_ = ~new_n7677_;
  assign new_n7699_ = new_n7701_ & new_n5722_;
  assign new_n7199_ = ~new_n9632_;
  assign new_n4562_ = ~new_n7699_;
  assign new_n7713_ = new_n7491_ & new_n7537_;
  assign new_n4563_ = ~new_n7713_;
  assign new_n7716_ = new_n7540_ & new_n7489_;
  assign new_n4564_ = ~new_n7716_;
  assign new_n7719_ = new_n7722_ & new_n7513_;
  assign new_n4565_ = ~new_n7719_;
  assign new_n7724_ = new_n7609_ | REG1_REG_15_;
  assign new_n4566_ = ~new_n7724_;
  assign new_n7730_ = new_n7732_ | REG1_REG_13_;
  assign new_n7200_ = ~new_n7790_;
  assign new_n4567_ = ~new_n7730_;
  assign new_n7742_ = new_n7492_ & new_n7537_;
  assign new_n4568_ = ~new_n7742_;
  assign new_n7745_ = new_n7540_ & new_n7490_;
  assign new_n4569_ = ~new_n7745_;
  assign new_n7748_ = new_n7493_ & new_n7513_;
  assign new_n4570_ = ~new_n7748_;
  assign new_n7751_ = new_n7463_ & new_n7353_;
  assign new_n4571_ = ~new_n7751_;
  assign new_n7755_ = new_n7357_ & new_n7455_;
  assign new_n7201_ = ~new_n9641_;
  assign new_n4572_ = ~new_n7755_;
  assign new_n7759_ = new_n7464_ & new_n7354_;
  assign new_n4573_ = ~new_n7759_;
  assign new_n7763_ = new_n7505_ & new_n7510_;
  assign new_n4574_ = ~new_n7763_;
  assign new_n7770_ = REG2_REG_31_ & new_n7568_;
  assign new_n4575_ = ~new_n7770_;
  assign new_n7773_ = new_n8115_ & new_n7775_;
  assign new_n4576_ = ~new_n7773_;
  assign new_n7778_ = REG2_REG_30_ & new_n7568_;
  assign new_n7202_ = ~new_n9741_;
  assign new_n4577_ = ~new_n7778_;
  assign new_n7780_ = new_n7781_ & new_n8115_;
  assign new_n4578_ = ~new_n7780_;
  assign new_n7795_ = new_n7799_ & new_n8115_;
  assign new_n4579_ = ~new_n7795_;
  assign new_n7804_ = new_n7807_ & new_n7558_;
  assign new_n4580_ = ~new_n7804_;
  assign new_n7812_ = new_n7561_ & new_n7816_;
  assign new_n4581_ = ~new_n7812_;
  assign new_n7817_ = new_n7772_ & new_n7004_;
  assign new_n7203_ = ~new_n9818_;
  assign new_n4582_ = ~new_n7817_;
  assign new_n7824_ = new_n7558_ & new_n7827_;
  assign new_n4583_ = ~new_n7824_;
  assign new_n7831_ = new_n7561_ & new_n7833_;
  assign new_n4584_ = ~new_n7831_;
  assign new_n7834_ = new_n7772_ & new_n7005_;
  assign new_n4585_ = ~new_n7834_;
  assign new_n7841_ = new_n7844_ & new_n7558_;
  assign new_n4586_ = ~new_n7841_;
  assign new_n7848_ = new_n7850_ & new_n7561_;
  assign new_n7204_ = ~new_n10000_;
  assign new_n4587_ = ~new_n7848_;
  assign new_n7851_ = new_n7772_ & new_n7006_;
  assign new_n4588_ = ~new_n7851_;
  assign new_n7858_ = new_n7861_ & new_n7558_;
  assign new_n4589_ = ~new_n7858_;
  assign new_n7865_ = new_n7561_ & new_n7867_;
  assign new_n4590_ = ~new_n7865_;
  assign new_n7868_ = new_n7772_ & new_n7007_;
  assign new_n4591_ = ~new_n7868_;
  assign new_n7875_ = new_n7878_ & new_n7558_;
  assign new_n7044_ = ~new_n8536_;
  assign new_n7205_ = ~new_n8585_;
  assign new_n4592_ = ~new_n7875_;
  assign new_n7882_ = new_n7884_ & new_n7561_;
  assign new_n4593_ = ~new_n7882_;
  assign new_n7885_ = new_n7772_ & new_n7009_;
  assign new_n4594_ = ~new_n7885_;
  assign new_n7892_ = new_n7895_ & new_n7558_;
  assign new_n4595_ = ~new_n7892_;
  assign new_n7899_ = new_n7561_ & new_n7901_;
  assign new_n4596_ = ~new_n7899_;
  assign new_n7902_ = new_n7772_ & new_n7011_;
  assign new_n7206_ = ~new_n11016_;
  assign new_n4597_ = ~new_n7902_;
  assign new_n7909_ = new_n7558_ & new_n7912_;
  assign new_n4598_ = ~new_n7909_;
  assign new_n7916_ = new_n7293_ & new_n7561_;
  assign new_n4599_ = ~new_n7916_;
  assign new_n7919_ = new_n7772_ & new_n7012_;
  assign new_n4600_ = ~new_n7919_;
  assign new_n7926_ = new_n7929_ & new_n7558_;
  assign new_n4601_ = ~new_n7926_;
  assign new_n7933_ = new_n7561_ & new_n7935_;
  assign new_n7733_ = new_n7350_ & new_n7510_;
  assign new_n4602_ = ~new_n7933_;
  assign new_n7936_ = new_n7772_ & new_n7013_;
  assign new_n4603_ = ~new_n7936_;
  assign new_n7943_ = new_n7946_ & new_n7558_;
  assign new_n4604_ = ~new_n7943_;
  assign new_n7950_ = new_n7952_ & new_n7561_;
  assign new_n4605_ = ~new_n7950_;
  assign new_n7953_ = new_n7772_ & new_n7014_;
  assign new_n4606_ = ~new_n7953_;
  assign new_n7960_ = new_n7963_ & new_n7558_;
  assign new_n7207_ = ~new_n7733_;
  assign new_n4607_ = ~new_n7960_;
  assign new_n7967_ = new_n7561_ & new_n7969_;
  assign new_n4608_ = ~new_n7967_;
  assign new_n7970_ = new_n7772_ & new_n7015_;
  assign new_n4609_ = ~new_n7970_;
  assign new_n7977_ = new_n7558_ & new_n7980_;
  assign new_n4610_ = ~new_n7977_;
  assign new_n7984_ = new_n7986_ & new_n7561_;
  assign new_n4611_ = ~new_n7984_;
  assign new_n7987_ = new_n7772_ & new_n7016_;
  assign new_n7208_ = ~new_n10603_;
  assign new_n4612_ = ~new_n7987_;
  assign new_n7994_ = new_n7997_ & new_n7558_;
  assign new_n4613_ = ~new_n7994_;
  assign new_n8001_ = new_n7561_ & new_n8003_;
  assign new_n4614_ = ~new_n8001_;
  assign new_n8004_ = new_n7772_ & new_n7017_;
  assign new_n4615_ = ~new_n8004_;
  assign new_n8011_ = new_n7558_ & new_n8014_;
  assign new_n4616_ = ~new_n8011_;
  assign new_n8018_ = new_n8020_ & new_n7561_;
  assign new_n11357_ = new_n11248_ & new_n7516_;
  assign new_n4617_ = ~new_n8018_;
  assign new_n8021_ = new_n7772_ & new_n7018_;
  assign new_n4618_ = ~new_n8021_;
  assign new_n8028_ = new_n7558_ & new_n8031_;
  assign new_n4619_ = ~new_n8028_;
  assign new_n8035_ = new_n7561_ & new_n8037_;
  assign new_n4620_ = ~new_n8035_;
  assign new_n8038_ = new_n7772_ & new_n7019_;
  assign new_n4621_ = ~new_n8038_;
  assign new_n8045_ = new_n7558_ & new_n8048_;
  assign new_n7209_ = ~new_n11357_;
  assign new_n4622_ = ~new_n8045_;
  assign new_n8052_ = new_n7294_ & new_n7561_;
  assign new_n4623_ = ~new_n8052_;
  assign new_n8055_ = new_n7772_ & new_n7021_;
  assign new_n4624_ = ~new_n8055_;
  assign new_n8062_ = new_n8065_ & new_n7558_;
  assign new_n4625_ = ~new_n8062_;
  assign new_n8069_ = new_n7561_ & new_n8071_;
  assign new_n4626_ = ~new_n8069_;
  assign new_n8072_ = new_n7772_ & new_n7023_;
  assign new_n11393_ = new_n11090_ & new_n7511_;
  assign new_n4627_ = ~new_n8072_;
  assign new_n8079_ = new_n8082_ & new_n7558_;
  assign new_n4628_ = ~new_n8079_;
  assign new_n8086_ = new_n8088_ & new_n7561_;
  assign new_n4629_ = ~new_n8086_;
  assign new_n8089_ = new_n7772_ & new_n7024_;
  assign new_n4630_ = ~new_n8089_;
  assign new_n8096_ = new_n7558_ & new_n8099_;
  assign new_n4631_ = ~new_n8096_;
  assign new_n8103_ = new_n7561_ & new_n8105_;
  assign new_n7210_ = ~new_n11393_;
  assign new_n4632_ = ~new_n8103_;
  assign new_n8106_ = new_n7772_ & new_n7025_;
  assign new_n4633_ = ~new_n8106_;
  assign new_n8113_ = new_n8118_ & new_n7558_;
  assign new_n4634_ = ~new_n8113_;
  assign new_n8122_ = new_n8124_ & new_n7561_;
  assign new_n4635_ = ~new_n8122_;
  assign new_n8125_ = new_n7772_ & new_n7026_;
  assign new_n4636_ = ~new_n8125_;
  assign new_n8132_ = new_n8135_ & new_n7558_;
  assign new_n8972_ = new_n8969_ & new_n7399_;
  assign new_n4637_ = ~new_n8132_;
  assign new_n8139_ = new_n7561_ & new_n8141_;
  assign new_n4638_ = ~new_n8139_;
  assign new_n8142_ = new_n7772_ & new_n7027_;
  assign new_n4639_ = ~new_n8142_;
  assign new_n8149_ = new_n7558_ & new_n8153_;
  assign new_n4640_ = ~new_n8149_;
  assign new_n8157_ = new_n8159_ & new_n7561_;
  assign new_n4641_ = ~new_n8157_;
  assign new_n8160_ = new_n7772_ & new_n7028_;
  assign new_n7045_ = ~new_n10531_;
  assign new_n7211_ = ~new_n8972_;
  assign new_n4642_ = ~new_n8160_;
  assign new_n8167_ = new_n8170_ & new_n7558_;
  assign new_n4643_ = ~new_n8167_;
  assign new_n8174_ = new_n7561_ & new_n8176_;
  assign new_n4644_ = ~new_n8174_;
  assign new_n8177_ = new_n7772_ & new_n7029_;
  assign new_n4645_ = ~new_n8177_;
  assign new_n8184_ = new_n7558_ & new_n8188_;
  assign new_n4646_ = ~new_n8184_;
  assign new_n8192_ = new_n7561_ & new_n8194_;
  assign new_n9121_ = new_n9126_ & new_n7520_;
  assign new_n4647_ = ~new_n8192_;
  assign new_n8195_ = new_n7772_ & new_n7030_;
  assign new_n4648_ = ~new_n8195_;
  assign new_n8202_ = new_n8205_ & new_n7558_;
  assign new_n4649_ = ~new_n8202_;
  assign new_n8209_ = new_n7561_ & new_n8211_;
  assign new_n4650_ = ~new_n8209_;
  assign new_n8212_ = new_n7772_ & new_n7031_;
  assign new_n4651_ = ~new_n8212_;
  assign new_n8219_ = new_n8222_ & new_n7561_;
  assign new_n7212_ = ~new_n9121_;
  assign new_n4652_ = ~new_n8219_;
  assign new_n8226_ = new_n7814_ & new_n9173_;
  assign new_n4653_ = ~new_n8226_;
  assign new_n8228_ = new_n7772_ & new_n7032_;
  assign new_n4654_ = ~new_n8228_;
  assign new_n8235_ = new_n7558_ & new_n8238_;
  assign new_n4655_ = ~new_n8235_;
  assign new_n8242_ = new_n7561_ & new_n8244_;
  assign new_n4656_ = ~new_n8242_;
  assign new_n8245_ = new_n7772_ & new_n7034_;
  assign new_n10801_ = REG3_REG_21_ & new_n10810_;
  assign new_n4657_ = ~new_n8245_;
  assign new_n8252_ = new_n8256_ & new_n7558_;
  assign new_n4658_ = ~new_n8252_;
  assign new_n8260_ = REG3_REG_2_ & new_n7561_;
  assign new_n4659_ = ~new_n8260_;
  assign new_n8263_ = new_n7772_ & new_n7035_;
  assign new_n4660_ = ~new_n8263_;
  assign new_n8270_ = new_n7558_ & new_n8273_;
  assign new_n4661_ = ~new_n8270_;
  assign new_n8277_ = REG3_REG_1_ & new_n7561_;
  assign new_n7213_ = ~new_n10801_;
  assign new_n4662_ = ~new_n8277_;
  assign new_n8279_ = new_n7772_ & new_n7036_;
  assign new_n4663_ = ~new_n8279_;
  assign new_n8299_ = new_n7568_ | new_n7701_;
  assign new_n4664_ = ~new_n8299_;
  assign new_n8296_ = new_n7558_ & new_n7411_;
  assign new_n4665_ = ~new_n8296_;
  assign new_n8410_ = new_n8406_ | new_n6697_;
  assign new_n4666_ = ~new_n8410_;
  assign new_n8430_ = new_n10635_ & new_n9290_;
  assign new_n10440_ = new_n7388_ & new_n10334_;
  assign new_n4667_ = ~new_n8430_;
  assign new_n8427_ = new_n8433_ & new_n8454_;
  assign new_n4668_ = ~new_n8427_;
  assign new_n8441_ = new_n8444_ & new_n7524_;
  assign new_n4669_ = ~new_n8441_;
  assign new_n8446_ = new_n7539_ & new_n7344_;
  assign new_n4670_ = ~new_n8446_;
  assign new_n8434_ = new_n7794_ & new_n8292_;
  assign new_n4671_ = ~new_n8434_;
  assign new_n8447_ = new_n7794_ & new_n8450_;
  assign new_n7214_ = ~new_n10440_;
  assign new_n4672_ = ~new_n8447_;
  assign new_n8452_ = new_n7367_ & new_n7519_;
  assign new_n4673_ = ~new_n8452_;
  assign new_n8464_ = new_n7807_ & new_n8292_;
  assign new_n4674_ = ~new_n8464_;
  assign new_n8476_ = new_n7807_ & new_n8450_;
  assign new_n4675_ = ~new_n8476_;
  assign new_n8497_ = new_n8498_ & new_n8503_;
  assign new_n4676_ = ~new_n8497_;
  assign new_n8499_ = new_n8502_ & new_n8503_;
  assign new_n7215_ = ~new_n10278_;
  assign new_n4677_ = ~new_n8499_;
  assign new_n8506_ = new_n8450_ & new_n7827_;
  assign new_n4678_ = ~new_n8506_;
  assign new_n8509_ = new_n6078_ & new_n7070_;
  assign new_n4679_ = ~new_n8509_;
  assign new_n8520_ = new_n7292_ | new_n7391_;
  assign new_n4680_ = ~new_n8520_;
  assign new_n8529_ = new_n7844_ & new_n8292_;
  assign new_n4681_ = ~new_n8529_;
  assign new_n8539_ = new_n7844_ & new_n8450_;
  assign new_n7216_ = ~new_n10402_;
  assign new_n4682_ = ~new_n8539_;
  assign new_n8561_ = new_n7861_ & new_n8292_;
  assign new_n4683_ = ~new_n8561_;
  assign new_n8567_ = new_n7861_ & new_n8450_;
  assign new_n4684_ = ~new_n8567_;
  assign new_n8580_ = new_n7878_ & new_n8292_;
  assign new_n4685_ = ~new_n8580_;
  assign new_n8589_ = new_n7878_ & new_n8450_;
  assign new_n4686_ = ~new_n8589_;
  assign new_n8594_ = new_n7358_ & new_n7538_;
  assign new_n7217_ = ~new_n8777_;
  assign new_n4687_ = ~new_n8594_;
  assign new_n8606_ = new_n7895_ & new_n8292_;
  assign new_n4688_ = ~new_n8606_;
  assign new_n8632_ = new_n7895_ & new_n8450_;
  assign new_n4689_ = ~new_n8632_;
  assign new_n8647_ = new_n7912_ & new_n8292_;
  assign new_n4690_ = ~new_n8647_;
  assign new_n8655_ = new_n8450_ & new_n7912_;
  assign new_n4691_ = ~new_n8655_;
  assign new_n8662_ = new_n8668_ & new_n7166_;
  assign new_n7024_ = ~new_n8091_;
  assign new_n7046_ = ~new_n11341_;
  assign new_n7218_ = ~new_n9078_;
  assign new_n4692_ = ~new_n8662_;
  assign new_n8682_ = new_n7929_ & new_n8292_;
  assign new_n4693_ = ~new_n8682_;
  assign new_n8688_ = new_n7929_ & new_n8450_;
  assign new_n4694_ = ~new_n8688_;
  assign new_n8691_ = new_n6087_ & new_n8685_;
  assign new_n4695_ = ~new_n8691_;
  assign new_n8695_ = new_n8698_ & new_n7167_;
  assign new_n4696_ = ~new_n8695_;
  assign new_n8706_ = new_n7946_ & new_n8292_;
  assign new_n7219_ = ~new_n9137_;
  assign new_n4697_ = ~new_n8706_;
  assign new_n8720_ = new_n7964_ | new_n7947_;
  assign new_n4698_ = ~new_n8720_;
  assign new_n8717_ = new_n7946_ & new_n8450_;
  assign new_n4699_ = ~new_n8717_;
  assign new_n8722_ = new_n8727_ & new_n8673_;
  assign new_n4700_ = ~new_n8722_;
  assign new_n8739_ = new_n7963_ & new_n8292_;
  assign new_n4701_ = ~new_n8739_;
  assign new_n8745_ = new_n7963_ & new_n8450_;
  assign new_n7220_ = ~new_n9971_;
  assign new_n4702_ = ~new_n8745_;
  assign new_n8758_ = new_n7980_ & new_n8292_;
  assign new_n4703_ = ~new_n8758_;
  assign new_n8768_ = new_n7981_ | new_n7998_;
  assign new_n4704_ = ~new_n8768_;
  assign new_n8765_ = new_n8450_ & new_n7980_;
  assign new_n4705_ = ~new_n8765_;
  assign new_n8785_ = new_n7997_ & new_n8292_;
  assign new_n4706_ = ~new_n8785_;
  assign new_n8792_ = new_n7997_ & new_n8450_;
  assign new_n7221_ = ~new_n10068_;
  assign new_n4707_ = ~new_n8792_;
  assign new_n8802_ = new_n7998_ & new_n8774_;
  assign new_n4708_ = ~new_n8802_;
  assign new_n8804_ = new_n7370_ & new_n7536_;
  assign new_n4709_ = ~new_n8804_;
  assign new_n8816_ = new_n6095_ & new_n7042_;
  assign new_n4710_ = ~new_n8816_;
  assign new_n8813_ = new_n8014_ & new_n8292_;
  assign new_n4711_ = ~new_n8813_;
  assign new_n8831_ = new_n8015_ | new_n8032_;
  assign new_n7222_ = ~new_n9596_;
  assign new_n4712_ = ~new_n8831_;
  assign new_n8828_ = new_n8450_ & new_n8014_;
  assign new_n4713_ = ~new_n8828_;
  assign new_n8836_ = new_n6097_ & new_n8841_;
  assign new_n4714_ = ~new_n8836_;
  assign new_n8850_ = new_n8031_ & new_n8292_;
  assign new_n4715_ = ~new_n8850_;
  assign new_n8860_ = new_n8450_ & new_n8031_;
  assign new_n4716_ = ~new_n8860_;
  assign new_n8877_ = new_n8048_ & new_n8292_;
  assign new_n7223_ = ~new_n8788_;
  assign new_n4717_ = ~new_n8877_;
  assign new_n8886_ = new_n8049_ | new_n8066_;
  assign new_n4718_ = ~new_n8886_;
  assign new_n8883_ = new_n8450_ & new_n8048_;
  assign new_n4719_ = ~new_n8883_;
  assign new_n8907_ = new_n8065_ & new_n8292_;
  assign new_n4720_ = ~new_n8907_;
  assign new_n8914_ = new_n8065_ & new_n8450_;
  assign new_n4721_ = ~new_n8914_;
  assign new_n8922_ = new_n7518_ & new_n7436_;
  assign new_n8789_ = new_n7523_ & new_n7409_;
  assign new_n4722_ = ~new_n8922_;
  assign new_n8926_ = new_n7247_ & new_n7518_;
  assign new_n4723_ = ~new_n8926_;
  assign new_n8936_ = new_n8082_ & new_n8292_;
  assign new_n4724_ = ~new_n8936_;
  assign new_n8948_ = new_n8100_ | new_n8083_;
  assign new_n4725_ = ~new_n8948_;
  assign new_n8945_ = new_n8082_ & new_n8450_;
  assign new_n4726_ = ~new_n8945_;
  assign new_n8963_ = new_n6104_ & new_n7043_;
  assign new_n7224_ = ~new_n8789_;
  assign new_n4727_ = ~new_n8963_;
  assign new_n8960_ = new_n8099_ & new_n8292_;
  assign new_n4728_ = ~new_n8960_;
  assign new_n8975_ = new_n8450_ & new_n8099_;
  assign new_n4729_ = ~new_n8975_;
  assign new_n8977_ = new_n7125_ & new_n5811_;
  assign new_n4730_ = ~new_n8977_;
  assign new_n8997_ = new_n8118_ & new_n8292_;
  assign new_n4731_ = ~new_n8997_;
  assign new_n9012_ = new_n8119_ | new_n8136_;
  assign new_n7225_ = ~new_n8761_;
  assign new_n4732_ = ~new_n9012_;
  assign new_n9009_ = new_n8118_ & new_n8450_;
  assign new_n4733_ = ~new_n9009_;
  assign new_n9019_ = new_n7535_ & new_n7433_;
  assign new_n4734_ = ~new_n9019_;
  assign new_n9023_ = new_n7250_ & new_n7535_;
  assign new_n4735_ = ~new_n9023_;
  assign new_n9033_ = new_n8135_ & new_n8292_;
  assign new_n4736_ = ~new_n9033_;
  assign new_n9039_ = new_n8135_ & new_n8450_;
  assign new_n7226_ = ~new_n8617_;
  assign new_n4737_ = ~new_n9039_;
  assign new_n9056_ = new_n6109_ & new_n7403_;
  assign new_n4738_ = ~new_n9056_;
  assign new_n9054_ = new_n9057_ & new_n5816_;
  assign new_n4739_ = ~new_n9054_;
  assign new_n9051_ = new_n8153_ & new_n8292_;
  assign new_n4740_ = ~new_n9051_;
  assign new_n9069_ = new_n8171_ | new_n8154_;
  assign new_n4741_ = ~new_n9069_;
  assign new_n9066_ = new_n8450_ & new_n8153_;
  assign new_n10704_ = new_n10119_ & STATE_REG;
  assign new_n9710_ = new_n10170_ & new_n10171_;
  assign new_n4742_ = ~new_n9066_;
  assign new_n9086_ = new_n8170_ & new_n8292_;
  assign new_n4743_ = ~new_n9086_;
  assign new_n9094_ = new_n8170_ & new_n8450_;
  assign new_n4744_ = ~new_n9094_;
  assign new_n9103_ = new_n8171_ & new_n9075_;
  assign new_n4745_ = ~new_n9103_;
  assign new_n9119_ = new_n7212_ & new_n7508_;
  assign new_n4746_ = ~new_n9119_;
  assign new_n9117_ = new_n9120_ & new_n5820_;
  assign new_n7227_ = ~new_n9710_;
  assign new_n4747_ = ~new_n9117_;
  assign new_n9114_ = new_n8188_ & new_n8292_;
  assign new_n4748_ = ~new_n9114_;
  assign new_n9132_ = new_n8206_ | new_n8189_;
  assign new_n4749_ = ~new_n9132_;
  assign new_n9129_ = new_n8450_ & new_n8188_;
  assign new_n4750_ = ~new_n9129_;
  assign new_n9140_ = new_n7533_ & new_n7421_;
  assign new_n4751_ = ~new_n9140_;
  assign new_n9149_ = new_n8205_ & new_n8292_;
  assign new_n7228_ = ~new_n9723_;
  assign new_n4752_ = ~new_n9149_;
  assign new_n9159_ = new_n8205_ & new_n8450_;
  assign new_n4753_ = ~new_n9159_;
  assign new_n9168_ = new_n8206_ & new_n9173_;
  assign new_n4754_ = ~new_n9168_;
  assign new_n9170_ = new_n7237_ & new_n7533_;
  assign new_n4755_ = ~new_n9170_;
  assign new_n9181_ = new_n8223_ & new_n8292_;
  assign new_n4756_ = ~new_n9181_;
  assign new_n9188_ = new_n8450_ & new_n8223_;
  assign new_n7229_ = ~new_n8869_;
  assign new_n4757_ = ~new_n9188_;
  assign new_n9193_ = new_n8239_ & new_n7363_;
  assign new_n4758_ = ~new_n9193_;
  assign new_n9204_ = new_n8238_ & new_n8292_;
  assign new_n4759_ = ~new_n9204_;
  assign new_n9211_ = new_n8450_ & new_n8238_;
  assign new_n4760_ = ~new_n9211_;
  assign new_n9213_ = new_n8257_ & new_n9216_;
  assign new_n4761_ = ~new_n9213_;
  assign new_n9224_ = new_n8256_ & new_n8292_;
  assign new_n7230_ = ~new_n10122_;
  assign new_n4762_ = ~new_n9224_;
  assign new_n9231_ = new_n8256_ & new_n8450_;
  assign new_n4763_ = ~new_n9231_;
  assign new_n9237_ = new_n9228_ & new_n7126_;
  assign new_n4764_ = ~new_n9237_;
  assign new_n9252_ = new_n8273_ & new_n8292_;
  assign new_n4765_ = ~new_n9252_;
  assign new_n9259_ = new_n8450_ & new_n8273_;
  assign new_n4766_ = ~new_n9259_;
  assign new_n9266_ = new_n6121_ & new_n7411_;
  assign new_n7231_ = ~new_n8454_;
  assign new_n4767_ = ~new_n9266_;
  assign new_n9286_ = new_n6124_ & new_n5828_;
  assign new_n4768_ = ~new_n9286_;
  assign new_n9308_ = new_n9314_ & new_n9305_;
  assign new_n4769_ = ~new_n9308_;
  assign new_n9317_ = new_n9311_ & IR_REG_29_;
  assign new_n4770_ = ~new_n9317_;
  assign new_n9324_ = new_n6128_ & new_n9329_;
  assign new_n4771_ = ~new_n9324_;
  assign new_n9332_ = new_n6129_ & new_n9338_;
  assign new_n7232_ = ~new_n8483_;
  assign new_n4772_ = ~new_n9332_;
  assign new_n9341_ = new_n9311_ & IR_REG_26_;
  assign new_n4773_ = ~new_n9341_;
  assign new_n9346_ = new_n9350_ & new_n9351_;
  assign new_n4774_ = ~new_n9346_;
  assign new_n9355_ = new_n6130_ & new_n9361_;
  assign new_n4775_ = ~new_n9355_;
  assign new_n9364_ = new_n9311_ & IR_REG_23_;
  assign new_n4776_ = ~new_n9364_;
  assign new_n9370_ = new_n6131_ & new_n9376_;
  assign new_n7233_ = ~new_n8596_;
  assign new_n4777_ = ~new_n9370_;
  assign new_n9379_ = new_n9311_ & IR_REG_21_;
  assign new_n4778_ = ~new_n9379_;
  assign new_n9385_ = new_n6132_ & new_n9391_;
  assign new_n4779_ = ~new_n9385_;
  assign new_n4780_ = ~new_n11152_;
  assign new_n9394_ = new_n9311_ & IR_REG_19_;
  assign new_n4781_ = ~new_n9394_;
  assign new_n9399_ = new_n6133_ & new_n9405_;
  assign new_n4782_ = ~new_n9399_;
  assign new_n7234_ = ~new_n8637_;
  assign new_n4783_ = ~new_n10680_;
  assign new_n9408_ = new_n9311_ & IR_REG_17_;
  assign new_n4784_ = ~new_n9408_;
  assign new_n9413_ = new_n6134_ & new_n9419_;
  assign new_n4785_ = ~new_n9413_;
  assign new_n9422_ = new_n9311_ & IR_REG_15_;
  assign new_n4786_ = ~new_n9422_;
  assign new_n9428_ = new_n6135_ & new_n9434_;
  assign new_n4787_ = ~new_n9428_;
  assign new_n9437_ = new_n9311_ & IR_REG_13_;
  assign new_n7235_ = ~new_n8805_;
  assign new_n4788_ = ~new_n9437_;
  assign new_n9443_ = new_n6136_ & new_n9449_;
  assign new_n4789_ = ~new_n9443_;
  assign new_n9452_ = new_n9311_ & IR_REG_11_;
  assign new_n4790_ = ~new_n9452_;
  assign new_n9458_ = new_n6137_ & new_n9464_;
  assign new_n4791_ = ~new_n9458_;
  assign new_n9467_ = new_n9311_ & IR_REG_9_;
  assign new_n4792_ = ~new_n9467_;
  assign new_n9473_ = new_n6138_ & new_n9478_;
  assign new_n7047_ = ~new_n10704_;
  assign new_n7236_ = ~new_n9106_;
  assign new_n4793_ = ~new_n9473_;
  assign new_n9481_ = new_n9311_ & IR_REG_7_;
  assign new_n4794_ = ~new_n9481_;
  assign new_n9488_ = new_n6139_ & new_n9494_;
  assign new_n4795_ = ~new_n9488_;
  assign new_n9497_ = new_n9311_ & IR_REG_5_;
  assign new_n4796_ = ~new_n9497_;
  assign new_n9502_ = new_n6140_ & new_n9508_;
  assign new_n4797_ = ~new_n9502_;
  assign new_n9511_ = new_n6141_ & new_n9516_;
  assign new_n7237_ = ~new_n9173_;
  assign new_n4798_ = ~new_n9511_;
  assign new_n9519_ = new_n9311_ & IR_REG_2_;
  assign new_n4799_ = ~new_n9519_;
  assign new_n9526_ = new_n6142_ & new_n9532_;
  assign new_n4800_ = ~new_n9526_;
  assign new_n9545_ = new_n9548_ & new_n9043_;
  assign new_n4801_ = ~new_n9545_;
  assign new_n9556_ = new_n9565_ & new_n10172_;
  assign new_n4802_ = ~new_n9556_;
  assign new_n9573_ = new_n9548_ & new_n8454_;
  assign new_n7238_ = ~new_n9171_;
  assign new_n4803_ = ~new_n9573_;
  assign new_n9577_ = new_n7828_ & new_n7556_;
  assign new_n4804_ = ~new_n9577_;
  assign new_n9587_ = new_n9548_ & new_n8841_;
  assign new_n4805_ = ~new_n9587_;
  assign new_n9591_ = new_n8049_ & new_n7556_;
  assign new_n4806_ = ~new_n9591_;
  assign new_n9602_ = new_n9548_ & new_n8521_;
  assign new_n4807_ = ~new_n9602_;
  assign new_n9606_ = new_n7896_ & new_n7556_;
  assign new_n7239_ = ~new_n8553_;
  assign new_n4808_ = ~new_n9606_;
  assign new_n9617_ = new_n9548_ & new_n8952_;
  assign new_n4809_ = ~new_n9617_;
  assign new_n9621_ = new_n8119_ & new_n7556_;
  assign new_n4810_ = ~new_n9621_;
  assign new_n9643_ = new_n9646_ & new_n7301_;
  assign new_n4811_ = ~new_n9643_;
  assign new_n9635_ = new_n8239_ & new_n7556_;
  assign new_n4812_ = ~new_n9635_;
  assign new_n9652_ = new_n9548_ & new_n8728_;
  assign new_n7240_ = ~new_n8552_;
  assign new_n4813_ = ~new_n9652_;
  assign new_n9656_ = new_n7964_ & new_n7556_;
  assign new_n4814_ = ~new_n9656_;
  assign new_n9667_ = new_n9548_ & new_n7815_;
  assign new_n4815_ = ~new_n9667_;
  assign new_n9678_ = new_n9681_ & new_n8454_;
  assign new_n4816_ = ~new_n9678_;
  assign new_n9682_ = new_n11114_ & new_n8454_;
  assign new_n4817_ = ~new_n9682_;
  assign new_n9690_ = new_n9681_ & new_n8483_;
  assign new_n7241_ = ~new_n8674_;
  assign new_n4818_ = ~new_n9690_;
  assign new_n9686_ = new_n9583_ & new_n7368_;
  assign new_n4819_ = ~new_n9686_;
  assign new_n9692_ = new_n9694_ & new_n7073_;
  assign new_n4820_ = ~new_n9692_;
  assign new_n9696_ = new_n11114_ & new_n8483_;
  assign new_n4821_ = ~new_n9696_;
  assign new_n9671_ = new_n7808_ & new_n7556_;
  assign new_n4822_ = ~new_n9671_;
  assign new_n9702_ = new_n9548_ & new_n9025_;
  assign new_n7242_ = ~new_n8728_;
  assign new_n4823_ = ~new_n9702_;
  assign new_n9706_ = new_n8154_ & new_n7556_;
  assign new_n4824_ = ~new_n9706_;
  assign new_n9715_ = new_n9548_ & new_n9216_;
  assign new_n4825_ = ~new_n9715_;
  assign new_n9719_ = REG3_REG_1_ & new_n9726_;
  assign new_n4826_ = ~new_n9719_;
  assign new_n9731_ = new_n9548_ & new_n8637_;
  assign new_n4827_ = ~new_n9731_;
  assign new_n9743_ = new_n7051_ & new_n7295_;
  assign new_n7243_ = ~new_n8729_;
  assign new_n4828_ = ~new_n9743_;
  assign new_n9753_ = new_n9548_ & new_n8927_;
  assign new_n4829_ = ~new_n9753_;
  assign new_n9757_ = new_n8083_ & new_n7556_;
  assign new_n4830_ = ~new_n9757_;
  assign new_n9767_ = new_n9548_ & new_n8553_;
  assign new_n4831_ = ~new_n9767_;
  assign new_n9771_ = new_n7862_ & new_n7556_;
  assign new_n4832_ = ~new_n9771_;
  assign new_n9781_ = new_n9548_ & new_n8774_;
  assign new_n7244_ = ~new_n8750_;
  assign new_n4833_ = ~new_n9781_;
  assign new_n9785_ = new_n8015_ & new_n7556_;
  assign new_n4834_ = ~new_n9785_;
  assign new_n9795_ = new_n9548_ & new_n9106_;
  assign new_n4835_ = ~new_n9795_;
  assign new_n9799_ = new_n8206_ & new_n7556_;
  assign new_n4836_ = ~new_n9799_;
  assign new_n9808_ = new_n9548_ & new_n8750_;
  assign new_n4837_ = ~new_n9808_;
  assign new_n9820_ = new_n7052_ & new_n7300_;
  assign new_n7245_ = ~new_n8841_;
  assign new_n4838_ = ~new_n9820_;
  assign new_n9828_ = new_n9548_ & new_n8552_;
  assign new_n4839_ = ~new_n9828_;
  assign new_n9832_ = new_n7879_ & new_n7556_;
  assign new_n4840_ = ~new_n9832_;
  assign new_n9843_ = new_n9548_ & new_n9173_;
  assign new_n4841_ = ~new_n9843_;
  assign new_n9847_ = new_n9849_ & new_n9554_;
  assign new_n4842_ = ~new_n9847_;
  assign new_n9858_ = new_n9548_ & new_n9024_;
  assign new_n7048_ = ~new_n8731_;
  assign new_n7246_ = ~new_n8927_;
  assign new_n4843_ = ~new_n9858_;
  assign new_n9862_ = new_n8136_ & new_n7556_;
  assign new_n4844_ = ~new_n9862_;
  assign new_n9871_ = new_n9548_ & new_n10442_;
  assign new_n4845_ = ~new_n9871_;
  assign new_n9874_ = new_n9235_ & new_n7556_;
  assign new_n4846_ = ~new_n9874_;
  assign new_n9880_ = new_n9548_ & new_n8674_;
  assign new_n4847_ = ~new_n9880_;
  assign new_n9884_ = new_n7947_ & new_n7556_;
  assign new_n7247_ = ~new_n8928_;
  assign new_n4848_ = ~new_n9884_;
  assign new_n9891_ = new_n9548_ & new_n8869_;
  assign new_n4849_ = ~new_n9891_;
  assign new_n9908_ = new_n7049_ & new_n7416_;
  assign new_n4850_ = ~new_n9908_;
  assign new_n9895_ = new_n8066_ & new_n7556_;
  assign new_n4851_ = ~new_n9895_;
  assign new_n9917_ = new_n9548_ & new_n8596_;
  assign new_n4852_ = ~new_n9917_;
  assign new_n9921_ = new_n7913_ & new_n7556_;
  assign new_n7248_ = ~new_n8952_;
  assign new_n4853_ = ~new_n9921_;
  assign new_n9932_ = new_n9548_ & new_n8928_;
  assign new_n4854_ = ~new_n9932_;
  assign new_n9941_ = new_n9946_ & new_n7400_;
  assign new_n4855_ = ~new_n9941_;
  assign new_n9936_ = new_n8100_ & new_n7556_;
  assign new_n4856_ = ~new_n9936_;
  assign new_n9951_ = new_n9548_ & new_n8262_;
  assign new_n4857_ = ~new_n9951_;
  assign new_n9955_ = REG3_REG_2_ & new_n9726_;
  assign new_n7249_ = ~new_n9024_;
  assign new_n4858_ = ~new_n9955_;
  assign new_n9962_ = new_n9548_ & new_n8729_;
  assign new_n4859_ = ~new_n9962_;
  assign new_n9966_ = new_n7981_ & new_n7556_;
  assign new_n4860_ = ~new_n9966_;
  assign new_n9977_ = new_n9548_ & new_n9075_;
  assign new_n4861_ = ~new_n9977_;
  assign new_n9981_ = new_n8189_ & new_n7556_;
  assign new_n4862_ = ~new_n9981_;
  assign new_n9991_ = new_n9548_ & new_n8483_;
  assign new_n7250_ = ~new_n9025_;
  assign new_n4863_ = ~new_n9991_;
  assign new_n10003_ = new_n9775_ & new_n7299_;
  assign new_n4864_ = ~new_n10003_;
  assign new_n10008_ = new_n11114_ & new_n8552_;
  assign new_n4865_ = ~new_n10008_;
  assign new_n10010_ = new_n9681_ & new_n8552_;
  assign new_n4866_ = ~new_n10010_;
  assign new_n10016_ = new_n9681_ & new_n8521_;
  assign new_n4867_ = ~new_n10016_;
  assign new_n10012_ = new_n7359_ & new_n7373_;
  assign new_n7251_ = ~new_n9043_;
  assign new_n4868_ = ~new_n10012_;
  assign new_n10018_ = new_n11114_ & new_n8521_;
  assign new_n4869_ = ~new_n10018_;
  assign new_n10024_ = new_n9681_ & new_n8596_;
  assign new_n4870_ = ~new_n10024_;
  assign new_n10020_ = new_n7360_ & new_n7374_;
  assign new_n4871_ = ~new_n10020_;
  assign new_n10026_ = new_n11114_ & new_n8596_;
  assign new_n4872_ = ~new_n10026_;
  assign new_n10036_ = new_n11114_ & new_n8674_;
  assign new_n7252_ = ~new_n7609_;
  assign new_n4873_ = ~new_n10036_;
  assign new_n10038_ = new_n9681_ & new_n8674_;
  assign new_n4874_ = ~new_n10038_;
  assign new_n10047_ = new_n11114_ & new_n8729_;
  assign new_n4875_ = ~new_n10047_;
  assign new_n10052_ = new_n9817_ & new_n7072_;
  assign new_n4876_ = ~new_n10052_;
  assign new_n10057_ = new_n11114_ & new_n8774_;
  assign new_n4877_ = ~new_n10057_;
  assign new_n10059_ = new_n9681_ & new_n8774_;
  assign new_n7253_ = ~new_n8969_;
  assign new_n4878_ = ~new_n10059_;
  assign new_n10072_ = new_n11114_ & new_n8805_;
  assign new_n4879_ = ~new_n10072_;
  assign new_n10074_ = new_n9681_ & new_n8805_;
  assign new_n4880_ = ~new_n10074_;
  assign new_n10051_ = new_n9970_ & new_n7375_;
  assign new_n4881_ = ~new_n10051_;
  assign new_n10077_ = new_n9681_ & new_n8750_;
  assign new_n4882_ = ~new_n10077_;
  assign new_n10079_ = new_n11114_ & new_n8750_;
  assign new_n7254_ = ~new_n9126_;
  assign new_n4883_ = ~new_n10079_;
  assign new_n10082_ = new_n9681_ & new_n8729_;
  assign new_n4884_ = ~new_n10082_;
  assign new_n10085_ = new_n11114_ & new_n8728_;
  assign new_n4885_ = ~new_n10085_;
  assign new_n10087_ = new_n9681_ & new_n8728_;
  assign new_n4886_ = ~new_n10087_;
  assign new_n10028_ = new_n9925_ & new_n7383_;
  assign new_n4887_ = ~new_n10028_;
  assign new_n10089_ = new_n11114_ & new_n8637_;
  assign new_n11129_ = new_n11145_ & new_n7296_;
  assign new_n4888_ = ~new_n10089_;
  assign new_n10092_ = new_n9681_ & new_n8637_;
  assign new_n4889_ = ~new_n10092_;
  assign new_n10098_ = new_n11114_ & new_n8553_;
  assign new_n4890_ = ~new_n10098_;
  assign new_n10100_ = new_n9681_ & new_n8553_;
  assign new_n4891_ = ~new_n10100_;
  assign new_n9995_ = new_n7845_ & new_n7556_;
  assign new_n4892_ = ~new_n9995_;
  assign new_n10105_ = new_n9548_ & new_n8805_;
  assign new_n7049_ = ~new_n9905_;
  assign new_n7255_ = ~new_n11129_;
  assign new_n4893_ = ~new_n10105_;
  assign new_n10112_ = new_n10116_ & STATE_REG;
  assign new_n4894_ = ~new_n10112_;
  assign new_n10133_ = new_n7314_ & new_n7258_;
  assign new_n4895_ = ~new_n10133_;
  assign new_n10131_ = new_n6145_ & new_n7443_;
  assign new_n4896_ = ~new_n10131_;
  assign new_n10141_ = new_n9681_ & new_n8841_;
  assign new_n4897_ = ~new_n10141_;
  assign new_n10143_ = new_n11114_ & new_n8841_;
  assign new_n9269_ = new_n9292_ & new_n7547_;
  assign new_n4898_ = ~new_n10143_;
  assign new_n10148_ = new_n10152_ & new_n5882_;
  assign new_n4899_ = ~new_n10148_;
  assign new_n10181_ = new_n11114_ & new_n9171_;
  assign new_n4900_ = ~new_n10181_;
  assign new_n10188_ = new_n11114_ & new_n8262_;
  assign new_n4901_ = ~new_n10188_;
  assign new_n10190_ = new_n9681_ & new_n8262_;
  assign new_n4902_ = ~new_n10190_;
  assign new_n10197_ = new_n10201_ & new_n7377_;
  assign new_n7256_ = ~new_n9269_;
  assign new_n4903_ = ~new_n10197_;
  assign new_n10203_ = new_n11114_ & new_n10442_;
  assign new_n4904_ = ~new_n10203_;
  assign new_n10205_ = new_n9681_ & new_n10442_;
  assign new_n4905_ = ~new_n10205_;
  assign new_n10211_ = new_n11114_ & new_n9216_;
  assign new_n4906_ = ~new_n10211_;
  assign new_n10213_ = new_n9681_ & new_n9216_;
  assign new_n4907_ = ~new_n10213_;
  assign new_n10216_ = new_n9681_ & new_n9171_;
  assign new_n7257_ = ~new_n9216_;
  assign new_n4908_ = ~new_n10216_;
  assign new_n10222_ = new_n9681_ & new_n9173_;
  assign new_n4909_ = ~new_n10222_;
  assign new_n10224_ = new_n11114_ & new_n9173_;
  assign new_n4910_ = ~new_n10224_;
  assign new_n10175_ = new_n7280_ & new_n5887_;
  assign new_n4911_ = ~new_n10175_;
  assign new_n10231_ = new_n11114_ & new_n9106_;
  assign new_n4912_ = ~new_n10231_;
  assign new_n10233_ = new_n9681_ & new_n9106_;
  assign new_n10135_ = new_n10324_ & new_n9282_;
  assign new_n4913_ = ~new_n10233_;
  assign new_n10236_ = new_n11114_ & new_n9075_;
  assign new_n4914_ = ~new_n10236_;
  assign new_n10238_ = new_n9681_ & new_n9075_;
  assign new_n4915_ = ~new_n10238_;
  assign new_n10244_ = new_n11114_ & new_n9043_;
  assign new_n4916_ = ~new_n10244_;
  assign new_n10246_ = new_n9681_ & new_n9043_;
  assign new_n4917_ = ~new_n10246_;
  assign new_n10249_ = new_n9681_ & new_n9025_;
  assign new_n7258_ = ~new_n10135_;
  assign new_n4918_ = ~new_n10249_;
  assign new_n10251_ = new_n11114_ & new_n9025_;
  assign new_n4919_ = ~new_n10251_;
  assign new_n10254_ = new_n11114_ & new_n9024_;
  assign new_n4920_ = ~new_n10254_;
  assign new_n10256_ = new_n9681_ & new_n9024_;
  assign new_n4921_ = ~new_n10256_;
  assign new_n10258_ = new_n11114_ & new_n8952_;
  assign new_n4922_ = ~new_n10258_;
  assign new_n10261_ = new_n9681_ & new_n8952_;
  assign new_n7259_ = ~new_n10432_;
  assign new_n4923_ = ~new_n10261_;
  assign new_n10264_ = new_n11114_ & new_n8927_;
  assign new_n4924_ = ~new_n10264_;
  assign new_n10266_ = new_n9681_ & new_n8927_;
  assign new_n4925_ = ~new_n10266_;
  assign new_n10269_ = new_n9681_ & new_n8928_;
  assign new_n4926_ = ~new_n10269_;
  assign new_n10272_ = new_n9681_ & new_n8869_;
  assign new_n4927_ = ~new_n10272_;
  assign new_n10274_ = new_n11114_ & new_n8869_;
  assign new_n10432_ = new_n8596_ & new_n7538_;
  assign new_n4928_ = ~new_n10274_;
  assign new_n10124_ = new_n8032_ & new_n7556_;
  assign new_n4929_ = ~new_n10124_;
  assign new_n10285_ = new_n9300_ & new_n5890_;
  assign new_n4930_ = ~new_n10285_;
  assign new_n10300_ = new_n9300_ & new_n5894_;
  assign new_n4931_ = ~new_n10300_;
  assign new_n10320_ = new_n10322_ & B_REG;
  assign new_n4932_ = ~new_n10320_;
  assign new_n10379_ = new_n6153_ & new_n10381_;
  assign new_n7260_ = ~new_n10319_;
  assign new_n4933_ = ~new_n10379_;
  assign new_n10392_ = new_n7472_ & new_n5913_;
  assign new_n4934_ = ~new_n10392_;
  assign new_n10400_ = new_n6155_ & new_n7459_;
  assign new_n4935_ = ~new_n10400_;
  assign new_n10386_ = new_n10410_ & new_n10389_;
  assign new_n4936_ = ~new_n10386_;
  assign new_n10330_ = new_n10422_ & new_n9292_;
  assign new_n4937_ = ~new_n10330_;
  assign new_n10428_ = new_n6293_ | new_n6705_;
  assign new_n7261_ = ~new_n11159_;
  assign new_n4938_ = ~new_n10428_;
  assign new_n10437_ = new_n6296_ | new_n6706_;
  assign new_n4939_ = ~new_n10437_;
  assign new_n10424_ = new_n6299_ | new_n6707_;
  assign new_n4940_ = ~new_n10424_;
  assign new_n10448_ = new_n6298_ | new_n10454_;
  assign new_n4941_ = ~new_n10448_;
  assign new_n10456_ = new_n6301_ | new_n10463_;
  assign new_n4942_ = ~new_n10456_;
  assign new_n10473_ = new_n6157_ & new_n7469_;
  assign new_n7050_ = ~new_n9567_;
  assign new_n7262_ = ~new_n11066_;
  assign new_n4943_ = ~new_n10473_;
  assign new_n10483_ = new_n6159_ & new_n5916_;
  assign new_n4944_ = ~new_n10483_;
  assign new_n10488_ = new_n8536_ & new_n7477_;
  assign new_n4945_ = ~new_n10488_;
  assign new_n10491_ = new_n10495_ & new_n7310_;
  assign new_n4946_ = ~new_n10491_;
  assign new_n10517_ = new_n7055_ & new_n7417_;
  assign new_n4947_ = ~new_n10517_;
  assign new_n10529_ = new_n10531_ & new_n5917_;
  assign new_n7263_ = ~new_n10138_;
  assign new_n4948_ = ~new_n10529_;
  assign new_n10555_ = new_n10556_ & new_n5922_;
  assign new_n4949_ = ~new_n10555_;
  assign new_n10575_ = new_n10361_ & new_n5925_;
  assign new_n4950_ = ~new_n10575_;
  assign new_n10579_ = new_n6165_ & new_n5927_;
  assign new_n4951_ = ~new_n10579_;
  assign new_n10588_ = new_n10635_ & new_n11036_;
  assign new_n4952_ = ~new_n10588_;
  assign new_n10591_ = new_n10635_ & new_n7511_;
  assign new_n7264_ = ~new_n10316_;
  assign new_n4953_ = ~new_n10591_;
  assign new_n10594_ = new_n7446_ & new_n10635_;
  assign new_n4954_ = ~new_n10594_;
  assign new_n10597_ = new_n10635_ & new_n11066_;
  assign new_n4955_ = ~new_n10597_;
  assign new_n10607_ = new_n11159_ & new_n10635_;
  assign new_n4956_ = ~new_n10607_;
  assign new_n10609_ = new_n10635_ & new_n7449_;
  assign new_n4957_ = ~new_n10609_;
  assign new_n10612_ = new_n7517_ & new_n10635_;
  assign new_n10316_ = new_n11460_ & new_n7313_;
  assign new_n4958_ = ~new_n10612_;
  assign new_n10615_ = new_n7516_ & new_n10635_;
  assign new_n4959_ = ~new_n10615_;
  assign new_n10618_ = new_n10635_ & new_n11179_;
  assign new_n4960_ = ~new_n10618_;
  assign new_n10534_ = new_n6306_ | new_n6716_;
  assign new_n4961_ = ~new_n10534_;
  assign new_n10622_ = new_n6166_ & new_n10334_;
  assign new_n4962_ = ~new_n10622_;
  assign new_n10639_ = new_n10432_ & new_n7522_;
  assign new_n7265_ = ~new_n8413_;
  assign new_n4963_ = ~new_n10639_;
  assign new_n10644_ = new_n10542_ & new_n5929_;
  assign new_n4964_ = ~new_n10644_;
  assign new_n10647_ = new_n10635_ & new_n7448_;
  assign new_n4965_ = ~new_n10647_;
  assign new_n10650_ = new_n7460_ & new_n10635_;
  assign new_n4966_ = ~new_n10650_;
  assign new_n10656_ = new_n7463_ & new_n10635_;
  assign new_n4967_ = ~new_n10656_;
  assign new_n10658_ = IR_REG_31_ & new_n5931_;
  assign new_n7266_ = ~new_n8117_;
  assign new_n4968_ = ~new_n10658_;
  assign new_n10661_ = new_n10635_ & new_n7513_;
  assign new_n4969_ = ~new_n10661_;
  assign new_n10665_ = new_n10667_ & IR_REG_31_;
  assign new_n4970_ = ~new_n10665_;
  assign new_n10669_ = new_n10635_ & new_n7510_;
  assign new_n4971_ = ~new_n10669_;
  assign new_n10671_ = new_n7464_ & new_n10635_;
  assign new_n4972_ = ~new_n10671_;
  assign new_n10673_ = IR_REG_31_ & new_n5932_;
  assign new_n7267_ = ~new_n8152_;
  assign new_n4973_ = ~new_n10673_;
  assign new_n10676_ = new_n7540_ & new_n10635_;
  assign new_n4974_ = ~new_n10676_;
  assign new_n10678_ = IR_REG_31_ & new_n10680_;
  assign new_n4975_ = ~new_n10678_;
  assign new_n10653_ = new_n6310_ | new_n6719_;
  assign new_n4976_ = ~new_n10653_;
  assign new_n10683_ = new_n10635_ & new_n7537_;
  assign new_n4977_ = ~new_n10683_;
  assign new_n10687_ = new_n6169_ & IR_REG_31_;
  assign new_n7268_ = ~new_n8187_;
  assign new_n4978_ = ~new_n10687_;
  assign new_n10690_ = new_n7545_ & new_n10635_;
  assign new_n4979_ = ~new_n10690_;
  assign new_n10692_ = new_n10635_ & new_n7455_;
  assign new_n4980_ = ~new_n10692_;
  assign new_n10695_ = new_n10697_ & IR_REG_31_;
  assign new_n4981_ = ~new_n10695_;
  assign new_n10710_ = REG2_REG_31_ & new_n7563_;
  assign new_n4982_ = ~new_n10710_;
  assign new_n10719_ = REG2_REG_30_ & new_n7563_;
  assign new_n7269_ = ~new_n10323_;
  assign new_n4983_ = ~new_n10719_;
  assign new_n10725_ = REG1_REG_29_ & new_n10709_;
  assign new_n4984_ = ~new_n10725_;
  assign new_n10727_ = REG0_REG_29_ & new_n7562_;
  assign new_n4985_ = ~new_n10727_;
  assign new_n10735_ = REG1_REG_28_ & new_n10709_;
  assign new_n4986_ = ~new_n10735_;
  assign new_n10737_ = REG0_REG_28_ & new_n7562_;
  assign new_n4987_ = ~new_n10737_;
  assign new_n10745_ = REG1_REG_27_ & new_n10709_;
  assign new_n10323_ = new_n11465_ & new_n7401_;
  assign new_n4988_ = ~new_n10745_;
  assign new_n10747_ = REG0_REG_27_ & new_n7562_;
  assign new_n4989_ = ~new_n10747_;
  assign new_n10753_ = REG1_REG_26_ & new_n10709_;
  assign new_n4990_ = ~new_n10753_;
  assign new_n10755_ = REG0_REG_26_ & new_n7562_;
  assign new_n4991_ = ~new_n10755_;
  assign new_n10766_ = REG1_REG_25_ & new_n10709_;
  assign new_n4992_ = ~new_n10766_;
  assign new_n10768_ = REG0_REG_25_ & new_n7562_;
  assign new_n7051_ = ~new_n9745_;
  assign new_n7270_ = ~new_n8698_;
  assign new_n4993_ = ~new_n10768_;
  assign new_n10774_ = REG1_REG_24_ & new_n10709_;
  assign new_n4994_ = ~new_n10774_;
  assign new_n10776_ = REG0_REG_24_ & new_n7562_;
  assign new_n4995_ = ~new_n10776_;
  assign new_n10787_ = REG1_REG_23_ & new_n10709_;
  assign new_n4996_ = ~new_n10787_;
  assign new_n10789_ = REG0_REG_23_ & new_n7562_;
  assign new_n4997_ = ~new_n10789_;
  assign new_n10795_ = REG1_REG_22_ & new_n10709_;
  assign new_n8698_ = new_n7964_ & new_n8729_;
  assign new_n4998_ = ~new_n10795_;
  assign new_n10797_ = REG0_REG_22_ & new_n7562_;
  assign new_n4999_ = ~new_n10797_;
  assign new_n10806_ = REG1_REG_21_ & new_n10709_;
  assign new_n5000_ = ~new_n10806_;
  assign new_n10808_ = REG0_REG_21_ & new_n7562_;
  assign new_n5001_ = ~new_n10808_;
  assign new_n10815_ = REG1_REG_20_ & new_n10709_;
  assign new_n5002_ = ~new_n10815_;
  assign new_n10817_ = REG0_REG_20_ & new_n7562_;
  assign new_n9625_ = new_n10163_ & new_n10164_;
  assign new_n5003_ = ~new_n10817_;
  assign new_n10827_ = new_n10709_ & REG1_REG_19_;
  assign new_n5004_ = ~new_n10827_;
  assign new_n10829_ = REG0_REG_19_ & new_n7562_;
  assign new_n5005_ = ~new_n10829_;
  assign new_n10835_ = new_n10709_ & REG1_REG_18_;
  assign new_n5006_ = ~new_n10835_;
  assign new_n10837_ = REG0_REG_18_ & new_n7562_;
  assign new_n5007_ = ~new_n10837_;
  assign new_n10848_ = new_n10709_ & REG1_REG_17_;
  assign new_n7271_ = ~new_n9625_;
  assign new_n5008_ = ~new_n10848_;
  assign new_n10850_ = REG0_REG_17_ & new_n7562_;
  assign new_n5009_ = ~new_n10850_;
  assign new_n10856_ = new_n10709_ & REG1_REG_16_;
  assign new_n5010_ = ~new_n10856_;
  assign new_n10858_ = REG0_REG_16_ & new_n7562_;
  assign new_n5011_ = ~new_n10858_;
  assign new_n10869_ = new_n10709_ & REG1_REG_15_;
  assign new_n5012_ = ~new_n10869_;
  assign new_n10871_ = REG0_REG_15_ & new_n7562_;
  assign new_n9484_ = new_n11432_ & new_n11431_;
  assign new_n5013_ = ~new_n10871_;
  assign new_n10877_ = new_n10709_ & REG1_REG_14_;
  assign new_n5014_ = ~new_n10877_;
  assign new_n10879_ = REG0_REG_14_ & new_n7562_;
  assign new_n5015_ = ~new_n10879_;
  assign new_n10889_ = new_n10709_ & REG1_REG_13_;
  assign new_n5016_ = ~new_n10889_;
  assign new_n10891_ = REG0_REG_13_ & new_n7562_;
  assign new_n5017_ = ~new_n10891_;
  assign new_n10897_ = new_n10709_ & REG1_REG_12_;
  assign new_n7272_ = ~new_n9484_;
  assign new_n5018_ = ~new_n10897_;
  assign new_n10899_ = REG0_REG_12_ & new_n7562_;
  assign new_n5019_ = ~new_n10899_;
  assign new_n10910_ = REG1_REG_11_ & new_n10709_;
  assign new_n5020_ = ~new_n10910_;
  assign new_n10912_ = REG0_REG_11_ & new_n7562_;
  assign new_n5021_ = ~new_n10912_;
  assign new_n10918_ = new_n10709_ & REG1_REG_10_;
  assign new_n5022_ = ~new_n10918_;
  assign new_n10920_ = REG0_REG_10_ & new_n7562_;
  assign new_n9790_ = new_n10062_ & new_n10063_;
  assign new_n5023_ = ~new_n10920_;
  assign new_n10931_ = new_n10709_ & REG1_REG_9_;
  assign new_n5024_ = ~new_n10931_;
  assign new_n10933_ = REG0_REG_9_ & new_n7562_;
  assign new_n5025_ = ~new_n10933_;
  assign new_n10939_ = new_n10709_ & REG1_REG_8_;
  assign new_n5026_ = ~new_n10939_;
  assign new_n10941_ = REG0_REG_8_ & new_n7562_;
  assign new_n5027_ = ~new_n10941_;
  assign new_n10952_ = new_n10709_ & REG1_REG_7_;
  assign new_n7273_ = ~new_n9790_;
  assign new_n5028_ = ~new_n10952_;
  assign new_n10954_ = REG0_REG_7_ & new_n7562_;
  assign new_n5029_ = ~new_n10954_;
  assign new_n10961_ = REG1_REG_6_ & new_n10709_;
  assign new_n5030_ = ~new_n10961_;
  assign new_n10963_ = REG0_REG_6_ & new_n7562_;
  assign new_n5031_ = ~new_n10963_;
  assign new_n10971_ = new_n10709_ & REG1_REG_5_;
  assign new_n5032_ = ~new_n10971_;
  assign new_n10973_ = REG0_REG_5_ & new_n7562_;
  assign new_n9903_ = new_n10149_ & new_n10150_;
  assign new_n5033_ = ~new_n10973_;
  assign new_n10979_ = new_n10709_ & REG1_REG_4_;
  assign new_n5034_ = ~new_n10979_;
  assign new_n10981_ = REG0_REG_4_ & new_n7562_;
  assign new_n5035_ = ~new_n10981_;
  assign new_n10988_ = new_n10709_ & REG1_REG_3_;
  assign new_n5036_ = ~new_n10988_;
  assign new_n10990_ = new_n10729_ & new_n8244_;
  assign new_n5037_ = ~new_n10990_;
  assign new_n10996_ = new_n10709_ & REG1_REG_2_;
  assign new_n7274_ = ~new_n9903_;
  assign new_n5038_ = ~new_n10996_;
  assign new_n10998_ = REG3_REG_2_ & new_n10729_;
  assign new_n5039_ = ~new_n10998_;
  assign new_n11004_ = REG1_REG_1_ & new_n10709_;
  assign new_n5040_ = ~new_n11004_;
  assign new_n11006_ = REG3_REG_1_ & new_n10729_;
  assign new_n5041_ = ~new_n11006_;
  assign new_n11012_ = REG3_REG_0_ & n1332;
  assign new_n5042_ = ~new_n11012_;
  assign new_n11026_ = REG3_REG_1_ & n1332;
  assign new_n7052_ = ~new_n9821_;
  assign new_n9002_ = new_n7453_ & new_n7399_;
  assign new_n5043_ = ~new_n11026_;
  assign new_n11030_ = new_n7580_ & new_n11037_;
  assign new_n5044_ = ~new_n11030_;
  assign new_n11044_ = new_n10596_ & new_n5967_;
  assign new_n5045_ = ~new_n11044_;
  assign new_n11059_ = ADDR_REG_2_ & new_n11294_;
  assign new_n5046_ = ~new_n11059_;
  assign new_n11064_ = new_n6204_ & new_n11066_;
  assign new_n5047_ = ~new_n11064_;
  assign new_n11084_ = new_n6206_ & new_n7511_;
  assign new_n7275_ = ~new_n9002_;
  assign new_n5048_ = ~new_n11084_;
  assign new_n11112_ = new_n11114_ & new_n10586_;
  assign new_n5049_ = ~new_n11112_;
  assign new_n11118_ = new_n7550_ & new_n7701_;
  assign new_n5050_ = ~new_n11118_;
  assign new_n11124_ = new_n9278_ | new_n9540_;
  assign new_n5051_ = ~new_n11124_;
  assign new_n11127_ = new_n7550_ | new_n7701_;
  assign new_n5052_ = ~new_n11127_;
  assign new_n11128_ = new_n7545_ | new_n7550_;
  assign new_n11397_ = new_n7483_ & new_n9508_;
  assign new_n5053_ = ~new_n11128_;
  assign new_n11122_ = new_n9681_ & new_n10586_;
  assign new_n5054_ = ~new_n11122_;
  assign new_n11134_ = new_n10709_ & REG1_REG_0_;
  assign new_n5055_ = ~new_n11134_;
  assign new_n11139_ = REG3_REG_0_ & new_n10729_;
  assign new_n5056_ = ~new_n11139_;
  assign new_n11141_ = IR_REG_31_ & new_n7162_;
  assign new_n5057_ = ~new_n11141_;
  assign new_n11144_ = new_n7550_ | new_n11129_;
  assign new_n7276_ = ~new_n11397_;
  assign new_n5058_ = ~new_n11144_;
  assign new_n11147_ = new_n6210_ & IR_REG_31_;
  assign new_n5059_ = ~new_n11147_;
  assign new_n11150_ = IR_REG_31_ & new_n11152_;
  assign new_n5060_ = ~new_n11150_;
  assign new_n11100_ = ADDR_REG_4_ & new_n11294_;
  assign new_n5061_ = ~new_n11100_;
  assign new_n11157_ = new_n11159_ & new_n5975_;
  assign new_n5062_ = ~new_n11157_;
  assign new_n11177_ = new_n6212_ & new_n11179_;
  assign new_n9777_ = new_n10004_ & new_n10005_;
  assign new_n5063_ = ~new_n11177_;
  assign new_n11198_ = new_n10614_ & new_n5980_;
  assign new_n5064_ = ~new_n11198_;
  assign new_n11217_ = new_n6215_ & new_n7449_;
  assign new_n5065_ = ~new_n11217_;
  assign new_n11236_ = new_n10617_ & new_n5986_;
  assign new_n5066_ = ~new_n11236_;
  assign new_n11255_ = new_n6218_ & new_n7448_;
  assign new_n5067_ = ~new_n11255_;
  assign new_n11274_ = new_n10652_ & new_n5992_;
  assign new_n7277_ = ~new_n9777_;
  assign new_n5068_ = ~new_n11274_;
  assign new_n11295_ = new_n6221_ & new_n7510_;
  assign new_n5069_ = ~new_n11295_;
  assign new_n11305_ = new_n11307_ & IR_REG_31_;
  assign new_n5070_ = ~new_n11305_;
  assign new_n11311_ = new_n7460_ & new_n7496_;
  assign new_n5071_ = ~new_n11311_;
  assign new_n11314_ = new_n7500_ & new_n7448_;
  assign new_n5072_ = ~new_n11314_;
  assign new_n11317_ = new_n7516_ & new_n7497_;
  assign new_n9744_ = new_n10041_ & new_n10042_;
  assign new_n5073_ = ~new_n11317_;
  assign new_n11320_ = new_n7501_ & new_n7449_;
  assign new_n5074_ = ~new_n11320_;
  assign new_n11323_ = new_n7517_ & new_n7498_;
  assign new_n5075_ = ~new_n11323_;
  assign new_n11326_ = new_n7502_ & new_n11179_;
  assign new_n5076_ = ~new_n11326_;
  assign new_n11329_ = new_n11159_ & new_n7494_;
  assign new_n5077_ = ~new_n11329_;
  assign new_n11332_ = new_n7503_ & new_n7511_;
  assign new_n7278_ = ~new_n9744_;
  assign new_n5078_ = ~new_n11332_;
  assign new_n11335_ = new_n7504_ & new_n11066_;
  assign new_n5079_ = ~new_n11335_;
  assign new_n11338_ = new_n7446_ & new_n7046_;
  assign new_n5080_ = ~new_n11338_;
  assign new_n11342_ = new_n7364_ & new_n11036_;
  assign new_n5081_ = ~new_n11342_;
  assign new_n11350_ = IR_REG_31_ & new_n5996_;
  assign new_n5082_ = ~new_n11350_;
  assign new_n11354_ = new_n11356_ | REG1_REG_10_;
  assign new_n9644_ = new_n10207_ & new_n10208_;
  assign new_n5083_ = ~new_n11354_;
  assign new_n11359_ = new_n6225_ & IR_REG_31_;
  assign new_n5084_ = ~new_n11359_;
  assign new_n11365_ = IR_REG_31_ & new_n5997_;
  assign new_n5085_ = ~new_n11365_;
  assign new_n11376_ = new_n6226_ & IR_REG_8_;
  assign new_n5086_ = ~new_n11376_;
  assign new_n11386_ = new_n6228_ & IR_REG_6_;
  assign new_n5087_ = ~new_n11386_;
  assign new_n11390_ = new_n11392_ | REG1_REG_5_;
  assign new_n7279_ = ~new_n9644_;
  assign new_n5088_ = ~new_n11390_;
  assign new_n11394_ = new_n9499_ & IR_REG_31_;
  assign new_n5089_ = ~new_n11394_;
  assign new_n11402_ = new_n6229_ & IR_REG_4_;
  assign new_n5090_ = ~new_n11402_;
  assign new_n11412_ = new_n6230_ & IR_REG_3_;
  assign new_n5091_ = ~new_n11412_;
  assign new_n11418_ = new_n7432_ & new_n11036_;
  assign new_n5092_ = ~new_n11418_;
  assign new_n11422_ = new_n6231_ & IR_REG_31_;
  assign new_n9154_ = new_n7520_ & new_n7508_;
  assign new_n9561_ = new_n10235_ & new_n10228_;
  assign new_n5093_ = ~new_n11422_;
  assign new_n11425_ = IR_REG_31_ & new_n5998_;
  assign new_n5094_ = ~new_n11425_;
  assign new_n11429_ = IR_REG_31_ & new_n5999_;
  assign new_n5095_ = ~new_n11429_;
  assign new_n11438_ = IR_REG_31_ & new_n6000_;
  assign new_n5096_ = ~new_n11438_;
  assign new_n11443_ = new_n6232_ & IR_REG_31_;
  assign new_n5097_ = ~new_n11443_;
  assign new_n11448_ = new_n6233_ & IR_REG_31_;
  assign new_n7280_ = ~new_n9561_;
  assign new_n5098_ = ~new_n11448_;
  assign new_n11452_ = new_n6234_ & IR_REG_31_;
  assign new_n5099_ = ~new_n11452_;
  assign new_n11436_ = new_n9540_ & new_n7450_;
  assign new_n5100_ = ~new_n11436_;
  assign new_n11433_ = new_n7056_ & new_n7047_;
  assign new_n5101_ = ~new_n11433_;
  assign new_n11456_ = IR_REG_31_ & new_n6001_;
  assign new_n5102_ = ~new_n11456_;
  assign new_n11455_ = new_n9540_ | n1332;
  assign new_n10465_ = new_n7445_ & new_n8952_;
  assign new_n5103_ = ~new_n11455_;
  assign new_n11462_ = new_n11464_ & IR_REG_31_;
  assign new_n5104_ = ~new_n11462_;
  assign new_n11466_ = new_n6235_ & IR_REG_31_;
  assign new_n5105_ = ~new_n11466_;
  assign new_n11469_ = new_n7150_ & IR_REG_31_;
  assign new_n5106_ = ~new_n11469_;
  assign new_n7573_ = ADDR_REG_13_ & new_n11294_;
  assign new_n5107_ = ~new_n7573_;
  assign new_n7575_ = new_n7464_ & new_n5707_;
  assign new_n7281_ = ~new_n10465_;
  assign new_n5108_ = ~new_n7575_;
  assign new_n7595_ = ADDR_REG_14_ & new_n11294_;
  assign new_n5109_ = ~new_n7595_;
  assign new_n7597_ = new_n7605_ & new_n5709_;
  assign new_n5110_ = ~new_n7597_;
  assign new_n7614_ = ADDR_REG_15_ & new_n11294_;
  assign new_n5111_ = ~new_n7614_;
  assign new_n7616_ = new_n7463_ & new_n5710_;
  assign new_n5112_ = ~new_n7616_;
  assign new_n7633_ = ADDR_REG_16_ & new_n11294_;
  assign new_n7282_ = ~new_n8840_;
  assign new_n5113_ = ~new_n7633_;
  assign new_n7635_ = new_n7646_ & new_n5712_;
  assign new_n5114_ = ~new_n7635_;
  assign new_n7648_ = new_n7586_ & new_n7649_;
  assign new_n5115_ = ~new_n7648_;
  assign new_n7654_ = ADDR_REG_17_ & new_n11294_;
  assign new_n5116_ = ~new_n7654_;
  assign new_n7656_ = new_n7540_ & new_n5714_;
  assign new_n5117_ = ~new_n7656_;
  assign new_n7676_ = ADDR_REG_18_ & new_n11294_;
  assign new_n11442_ = new_n7466_ & new_n9376_;
  assign new_n5118_ = ~new_n7676_;
  assign new_n7678_ = new_n7689_ & new_n5718_;
  assign new_n5119_ = ~new_n7678_;
  assign new_n7692_ = new_n7586_ & new_n7693_;
  assign new_n5120_ = ~new_n7692_;
  assign new_n7698_ = ADDR_REG_19_ & new_n11294_;
  assign new_n5121_ = ~new_n7698_;
  assign new_n7700_ = new_n7545_ & new_n5720_;
  assign new_n5122_ = ~new_n7700_;
  assign new_n7714_ = new_n7715_ & new_n7684_;
  assign new_n7283_ = ~new_n11442_;
  assign new_n5123_ = ~new_n7714_;
  assign new_n7717_ = new_n7718_ & new_n7669_;
  assign new_n5124_ = ~new_n7717_;
  assign new_n7720_ = new_n6012_ & new_n7640_;
  assign new_n5125_ = ~new_n7720_;
  assign new_n7723_ = new_n7617_ & new_n7093_;
  assign new_n5126_ = ~new_n7723_;
  assign new_n7726_ = new_n7119_ & new_n7252_;
  assign new_n5127_ = ~new_n7726_;
  assign new_n7727_ = new_n7120_ & new_n7304_;
  assign new_n10660_ = new_n7397_ & new_n9434_;
  assign new_n5128_ = ~new_n7727_;
  assign new_n7743_ = new_n7744_ & new_n7688_;
  assign new_n5129_ = ~new_n7743_;
  assign new_n7746_ = new_n7747_ & new_n7672_;
  assign new_n5130_ = ~new_n7746_;
  assign new_n7749_ = new_n7750_ & new_n7644_;
  assign new_n5131_ = ~new_n7749_;
  assign new_n7752_ = new_n7753_ & new_n7754_;
  assign new_n5132_ = ~new_n7752_;
  assign new_n7756_ = new_n7757_ & new_n7758_;
  assign new_n7284_ = ~new_n10660_;
  assign new_n5133_ = ~new_n7756_;
  assign new_n7760_ = new_n7761_ & new_n7762_;
  assign new_n5134_ = ~new_n7760_;
  assign new_n7764_ = new_n7765_ & new_n7766_;
  assign new_n5135_ = ~new_n7764_;
  assign new_n7771_ = new_n7809_ & new_n8404_;
  assign new_n5136_ = ~new_n7771_;
  assign new_n7779_ = new_n8416_ & new_n7809_;
  assign new_n5137_ = ~new_n7779_;
  assign new_n7787_ = new_n8415_ & new_n7809_;
  assign new_n10675_ = new_n7398_ & new_n9449_;
  assign new_n5138_ = ~new_n7787_;
  assign new_n7792_ = new_n7558_ & new_n7794_;
  assign new_n5139_ = ~new_n7792_;
  assign new_n7805_ = new_n7806_ & new_n8115_;
  assign new_n5140_ = ~new_n7805_;
  assign new_n7813_ = new_n7814_ & new_n7815_;
  assign new_n5141_ = ~new_n7813_;
  assign new_n7818_ = REG2_REG_28_ & new_n7568_;
  assign new_n5142_ = ~new_n7818_;
  assign new_n7825_ = new_n7826_ & new_n8115_;
  assign new_n7053_ = ~new_n9154_;
  assign new_n7285_ = ~new_n10675_;
  assign new_n5143_ = ~new_n7825_;
  assign new_n7832_ = new_n7814_ & new_n8454_;
  assign new_n5144_ = ~new_n7832_;
  assign new_n7835_ = REG2_REG_27_ & new_n7568_;
  assign new_n5145_ = ~new_n7835_;
  assign new_n7842_ = new_n7843_ & new_n8115_;
  assign new_n5146_ = ~new_n7842_;
  assign new_n7849_ = new_n7814_ & new_n8483_;
  assign new_n5147_ = ~new_n7849_;
  assign new_n7852_ = REG2_REG_26_ & new_n7568_;
  assign new_n11352_ = new_n7467_ & new_n9464_;
  assign new_n5148_ = ~new_n7852_;
  assign new_n7859_ = new_n7860_ & new_n8115_;
  assign new_n5149_ = ~new_n7859_;
  assign new_n7866_ = new_n7814_ & new_n8553_;
  assign new_n5150_ = ~new_n7866_;
  assign new_n7869_ = REG2_REG_25_ & new_n7568_;
  assign new_n5151_ = ~new_n7869_;
  assign new_n7876_ = new_n7877_ & new_n8115_;
  assign new_n5152_ = ~new_n7876_;
  assign new_n7883_ = new_n7814_ & new_n8552_;
  assign new_n7286_ = ~new_n11352_;
  assign new_n5153_ = ~new_n7883_;
  assign new_n7886_ = REG2_REG_24_ & new_n7568_;
  assign new_n5154_ = ~new_n7886_;
  assign new_n7893_ = new_n7894_ & new_n8115_;
  assign new_n5155_ = ~new_n7893_;
  assign new_n7900_ = new_n7814_ & new_n8521_;
  assign new_n5156_ = ~new_n7900_;
  assign new_n7903_ = REG2_REG_23_ & new_n7568_;
  assign new_n5157_ = ~new_n7903_;
  assign new_n7910_ = new_n7911_ & new_n8115_;
  assign new_n11368_ = new_n9484_ & new_n9478_;
  assign new_n5158_ = ~new_n7910_;
  assign new_n7917_ = new_n7814_ & new_n8596_;
  assign new_n5159_ = ~new_n7917_;
  assign new_n7920_ = REG2_REG_22_ & new_n7568_;
  assign new_n5160_ = ~new_n7920_;
  assign new_n7927_ = new_n7928_ & new_n8115_;
  assign new_n5161_ = ~new_n7927_;
  assign new_n7934_ = new_n7814_ & new_n8637_;
  assign new_n5162_ = ~new_n7934_;
  assign new_n7937_ = REG2_REG_21_ & new_n7568_;
  assign new_n7287_ = ~new_n11368_;
  assign new_n5163_ = ~new_n7937_;
  assign new_n7944_ = new_n7945_ & new_n8115_;
  assign new_n5164_ = ~new_n7944_;
  assign new_n7951_ = new_n7814_ & new_n8674_;
  assign new_n5165_ = ~new_n7951_;
  assign new_n7954_ = REG2_REG_20_ & new_n7568_;
  assign new_n5166_ = ~new_n7954_;
  assign new_n7961_ = new_n8115_ & new_n7962_;
  assign new_n5167_ = ~new_n7961_;
  assign new_n7968_ = new_n7814_ & new_n8728_;
  assign new_n9241_ = new_n8274_ & new_n10442_;
  assign new_n5168_ = ~new_n7968_;
  assign new_n7971_ = REG2_REG_19_ & new_n7568_;
  assign new_n5169_ = ~new_n7971_;
  assign new_n7978_ = new_n7979_ & new_n8115_;
  assign new_n5170_ = ~new_n7978_;
  assign new_n7985_ = new_n7814_ & new_n8729_;
  assign new_n5171_ = ~new_n7985_;
  assign new_n7988_ = REG2_REG_18_ & new_n7568_;
  assign new_n5172_ = ~new_n7988_;
  assign new_n7995_ = new_n8115_ & new_n7996_;
  assign new_n7288_ = ~new_n9241_;
  assign new_n5173_ = ~new_n7995_;
  assign new_n8002_ = new_n7814_ & new_n8750_;
  assign new_n5174_ = ~new_n8002_;
  assign new_n8005_ = REG2_REG_17_ & new_n7568_;
  assign new_n5175_ = ~new_n8005_;
  assign new_n8012_ = new_n8013_ & new_n8115_;
  assign new_n5176_ = ~new_n8012_;
  assign new_n8019_ = new_n7814_ & new_n8774_;
  assign new_n5177_ = ~new_n8019_;
  assign new_n8022_ = REG2_REG_16_ & new_n7568_;
  assign new_n7289_ = ~new_n10464_;
  assign new_n5178_ = ~new_n8022_;
  assign new_n8029_ = new_n8115_ & new_n8030_;
  assign new_n5179_ = ~new_n8029_;
  assign new_n8036_ = new_n7814_ & new_n8805_;
  assign new_n5180_ = ~new_n8036_;
  assign new_n8039_ = REG2_REG_15_ & new_n7568_;
  assign new_n5181_ = ~new_n8039_;
  assign new_n8046_ = new_n8047_ & new_n8115_;
  assign new_n5182_ = ~new_n8046_;
  assign new_n8053_ = new_n7814_ & new_n8841_;
  assign new_n9564_ = new_n10218_ & new_n10219_;
  assign new_n5183_ = ~new_n8053_;
  assign new_n8056_ = REG2_REG_14_ & new_n7568_;
  assign new_n5184_ = ~new_n8056_;
  assign new_n8063_ = new_n8115_ & new_n8064_;
  assign new_n5185_ = ~new_n8063_;
  assign new_n8070_ = new_n7814_ & new_n8869_;
  assign new_n5186_ = ~new_n8070_;
  assign new_n8073_ = REG2_REG_13_ & new_n7568_;
  assign new_n5187_ = ~new_n8073_;
  assign new_n8080_ = new_n8081_ & new_n8115_;
  assign new_n7290_ = ~new_n9564_;
  assign new_n5188_ = ~new_n8080_;
  assign new_n8087_ = new_n7814_ & new_n8927_;
  assign new_n5189_ = ~new_n8087_;
  assign new_n8090_ = REG2_REG_12_ & new_n7568_;
  assign new_n5190_ = ~new_n8090_;
  assign new_n8097_ = new_n8115_ & new_n8098_;
  assign new_n5191_ = ~new_n8097_;
  assign new_n8104_ = new_n7814_ & new_n8928_;
  assign new_n5192_ = ~new_n8104_;
  assign new_n8107_ = REG2_REG_11_ & new_n7568_;
  assign new_n7025_ = ~new_n8108_;
  assign new_n7054_ = ~new_n10378_;
  assign new_n7291_ = ~new_n9626_;
  assign new_n5193_ = ~new_n8107_;
  assign new_n8123_ = new_n7814_ & new_n8952_;
  assign new_n5194_ = ~new_n8123_;
  assign new_n8126_ = REG2_REG_10_ & new_n7568_;
  assign new_n5195_ = ~new_n8126_;
  assign new_n8133_ = new_n8115_ & new_n8134_;
  assign new_n5196_ = ~new_n8133_;
  assign new_n8140_ = new_n7814_ & new_n9024_;
  assign new_n5197_ = ~new_n8140_;
  assign new_n8143_ = REG2_REG_9_ & new_n7568_;
  assign new_n7292_ = ~new_n8512_;
  assign new_n5198_ = ~new_n8143_;
  assign new_n8158_ = new_n7814_ & new_n9025_;
  assign new_n5199_ = ~new_n8158_;
  assign new_n8161_ = REG2_REG_8_ & new_n7568_;
  assign new_n5200_ = ~new_n8161_;
  assign new_n8168_ = new_n8115_ & new_n8169_;
  assign new_n5201_ = ~new_n8168_;
  assign new_n8175_ = new_n7814_ & new_n9043_;
  assign new_n5202_ = ~new_n8175_;
  assign new_n8178_ = REG2_REG_7_ & new_n7568_;
  assign new_n7918_ = new_n10799_ | new_n7439_;
  assign new_n5203_ = ~new_n8178_;
  assign new_n8193_ = new_n7814_ & new_n9075_;
  assign new_n5204_ = ~new_n8193_;
  assign new_n8196_ = REG2_REG_6_ & new_n7568_;
  assign new_n5205_ = ~new_n8196_;
  assign new_n8203_ = new_n8115_ & new_n8204_;
  assign new_n5206_ = ~new_n8203_;
  assign new_n8210_ = new_n7814_ & new_n9106_;
  assign new_n5207_ = ~new_n8210_;
  assign new_n8213_ = REG2_REG_5_ & new_n7568_;
  assign new_n7293_ = ~new_n7918_;
  assign new_n5208_ = ~new_n8213_;
  assign new_n8227_ = new_n9172_ & new_n7809_;
  assign new_n5209_ = ~new_n8227_;
  assign new_n8229_ = REG2_REG_4_ & new_n7568_;
  assign new_n5210_ = ~new_n8229_;
  assign new_n8236_ = new_n8115_ & new_n8237_;
  assign new_n5211_ = ~new_n8236_;
  assign new_n8243_ = new_n7814_ & new_n9171_;
  assign new_n5212_ = ~new_n8243_;
  assign new_n8246_ = REG2_REG_3_ & new_n7568_;
  assign new_n7294_ = ~new_n8054_;
  assign new_n5213_ = ~new_n8246_;
  assign new_n8261_ = new_n7814_ & new_n8262_;
  assign new_n5214_ = ~new_n8261_;
  assign new_n8264_ = REG2_REG_2_ & new_n7568_;
  assign new_n5215_ = ~new_n8264_;
  assign new_n8271_ = new_n8115_ & new_n8272_;
  assign new_n5216_ = ~new_n8271_;
  assign new_n8278_ = new_n7814_ & new_n9216_;
  assign new_n5217_ = ~new_n8278_;
  assign new_n8280_ = REG2_REG_1_ & new_n7568_;
  assign new_n7295_ = ~new_n9746_;
  assign new_n5218_ = ~new_n8280_;
  assign new_n8285_ = REG3_REG_0_ & new_n7561_;
  assign new_n5219_ = ~new_n8285_;
  assign new_n8294_ = new_n7814_ & new_n10442_;
  assign new_n5220_ = ~new_n8294_;
  assign new_n8298_ = new_n7544_ & new_n7559_;
  assign new_n5221_ = ~new_n8298_;
  assign new_n8403_ = new_n9269_ & new_n8404_;
  assign new_n5222_ = ~new_n8403_;
  assign new_n8411_ = new_n8416_ & new_n9269_;
  assign new_n11146_ = new_n7527_ & new_n9391_;
  assign new_n5223_ = ~new_n8411_;
  assign new_n8417_ = new_n8449_ & new_n7461_;
  assign new_n5224_ = ~new_n8417_;
  assign new_n8424_ = new_n8415_ & new_n9269_;
  assign new_n5225_ = ~new_n8424_;
  assign new_n8428_ = new_n7480_ & new_n7122_;
  assign new_n5226_ = ~new_n8428_;
  assign new_n8431_ = new_n8295_ & new_n8432_;
  assign new_n5227_ = ~new_n8431_;
  assign new_n8435_ = new_n6075_ & new_n7560_;
  assign new_n7296_ = ~new_n11146_;
  assign new_n5228_ = ~new_n8435_;
  assign new_n8448_ = new_n7799_ & new_n8413_;
  assign new_n5229_ = ~new_n8448_;
  assign new_n8453_ = new_n7231_ & new_n8455_;
  assign new_n5230_ = ~new_n8453_;
  assign new_n8461_ = new_n7808_ & new_n9269_;
  assign new_n5231_ = ~new_n8461_;
  assign new_n8463_ = new_n8433_ & new_n8483_;
  assign new_n5232_ = ~new_n8463_;
  assign new_n8469_ = new_n8470_ & new_n7435_;
  assign new_n9321_ = new_n11447_ & new_n9329_;
  assign new_n5233_ = ~new_n8469_;
  assign new_n8475_ = new_n8295_ & new_n7815_;
  assign new_n5234_ = ~new_n8475_;
  assign new_n8480_ = new_n8508_ & new_n7457_;
  assign new_n5235_ = ~new_n8480_;
  assign new_n8482_ = new_n7232_ & new_n5788_;
  assign new_n5236_ = ~new_n8482_;
  assign new_n8490_ = new_n7828_ & new_n9269_;
  assign new_n5237_ = ~new_n8490_;
  assign new_n8492_ = new_n8433_ & new_n8553_;
  assign new_n7297_ = ~new_n9321_;
  assign new_n5238_ = ~new_n8492_;
  assign new_n8500_ = new_n8501_ & new_n7514_;
  assign new_n5239_ = ~new_n8500_;
  assign new_n8505_ = new_n8295_ & new_n8454_;
  assign new_n5240_ = ~new_n8505_;
  assign new_n8510_ = new_n8511_ & new_n8512_;
  assign new_n5241_ = ~new_n8510_;
  assign new_n8526_ = new_n7845_ & new_n9269_;
  assign new_n5242_ = ~new_n8526_;
  assign new_n8528_ = new_n8433_ & new_n8552_;
  assign new_n10525_ = new_n7471_ & new_n7387_;
  assign new_n8517_ = new_n7862_ & new_n8552_;
  assign new_n5243_ = ~new_n8528_;
  assign new_n8534_ = new_n7487_ & new_n7044_;
  assign new_n5244_ = ~new_n8534_;
  assign new_n8538_ = new_n8295_ & new_n8483_;
  assign new_n5245_ = ~new_n8538_;
  assign new_n8543_ = new_n8569_ & new_n7512_;
  assign new_n5246_ = ~new_n8543_;
  assign new_n8550_ = new_n7298_ & new_n7008_;
  assign new_n5247_ = ~new_n8550_;
  assign new_n8558_ = new_n7862_ & new_n9269_;
  assign new_n7298_ = ~new_n8517_;
  assign new_n5248_ = ~new_n8558_;
  assign new_n8560_ = new_n8433_ & new_n8521_;
  assign new_n5249_ = ~new_n8560_;
  assign new_n8566_ = new_n8295_ & new_n8553_;
  assign new_n5250_ = ~new_n8566_;
  assign new_n8570_ = new_n6081_ & new_n7010_;
  assign new_n5251_ = ~new_n8570_;
  assign new_n8577_ = new_n7879_ & new_n9269_;
  assign new_n5252_ = ~new_n8577_;
  assign new_n8579_ = new_n8433_ & new_n8596_;
  assign new_n7299_ = ~new_n9776_;
  assign new_n5253_ = ~new_n8579_;
  assign new_n8588_ = new_n8295_ & new_n8552_;
  assign new_n5254_ = ~new_n8588_;
  assign new_n8593_ = new_n8634_ & new_n7538_;
  assign new_n5255_ = ~new_n8593_;
  assign new_n8595_ = new_n7233_ & new_n8597_;
  assign new_n5256_ = ~new_n8595_;
  assign new_n8603_ = new_n7896_ & new_n9269_;
  assign new_n5257_ = ~new_n8603_;
  assign new_n8605_ = new_n8433_ & new_n8637_;
  assign new_n7300_ = ~new_n9789_;
  assign new_n5258_ = ~new_n8605_;
  assign new_n8612_ = new_n6084_ & new_n7434_;
  assign new_n5259_ = ~new_n8612_;
  assign new_n8616_ = new_n7226_ & new_n7530_;
  assign new_n5260_ = ~new_n8616_;
  assign new_n8622_ = new_n7526_ & new_n7310_;
  assign new_n5261_ = ~new_n8622_;
  assign new_n8626_ = new_n8627_ & new_n7526_;
  assign new_n5262_ = ~new_n8626_;
  assign new_n8631_ = new_n8295_ & new_n8521_;
  assign new_n7301_ = ~new_n9645_;
  assign new_n5263_ = ~new_n8631_;
  assign new_n8636_ = new_n7234_ & new_n5794_;
  assign new_n5264_ = ~new_n8636_;
  assign new_n8644_ = new_n7913_ & new_n9269_;
  assign new_n5265_ = ~new_n8644_;
  assign new_n8646_ = new_n8433_ & new_n8674_;
  assign new_n5266_ = ~new_n8646_;
  assign new_n8651_ = new_n8652_ & new_n7526_;
  assign new_n5267_ = ~new_n8651_;
  assign new_n8654_ = new_n8295_ & new_n8596_;
  assign new_n7302_ = ~new_n10460_;
  assign new_n5268_ = ~new_n8654_;
  assign new_n8659_ = new_n8690_ & new_n7509_;
  assign new_n5269_ = ~new_n8659_;
  assign new_n8661_ = new_n7930_ & new_n8674_;
  assign new_n5270_ = ~new_n8661_;
  assign new_n8679_ = new_n7930_ & new_n9269_;
  assign new_n5271_ = ~new_n8679_;
  assign new_n8681_ = new_n8433_ & new_n8728_;
  assign new_n5272_ = ~new_n8681_;
  assign new_n8687_ = new_n8295_ & new_n8637_;
  assign new_n7303_ = ~new_n10602_;
  assign new_n5273_ = ~new_n8687_;
  assign new_n8703_ = new_n7947_ & new_n9269_;
  assign new_n5274_ = ~new_n8703_;
  assign new_n8705_ = new_n8433_ & new_n8729_;
  assign new_n5275_ = ~new_n8705_;
  assign new_n8712_ = new_n7484_ & new_n7365_;
  assign new_n5276_ = ~new_n8712_;
  assign new_n8716_ = new_n8295_ & new_n8674_;
  assign new_n5277_ = ~new_n8716_;
  assign new_n8721_ = new_n8747_ & new_n7438_;
  assign new_n7590_ = new_n7735_ & REG1_REG_13_;
  assign new_n5278_ = ~new_n8721_;
  assign new_n8736_ = new_n7964_ & new_n9269_;
  assign new_n5279_ = ~new_n8736_;
  assign new_n8738_ = new_n8433_ & new_n8750_;
  assign new_n5280_ = ~new_n8738_;
  assign new_n8744_ = new_n8295_ & new_n8728_;
  assign new_n5281_ = ~new_n8744_;
  assign new_n8748_ = new_n8667_ & new_n5799_;
  assign new_n5282_ = ~new_n8748_;
  assign new_n8755_ = new_n7981_ & new_n9269_;
  assign new_n7304_ = ~new_n7590_;
  assign new_n5283_ = ~new_n8755_;
  assign new_n8757_ = new_n8433_ & new_n8774_;
  assign new_n5284_ = ~new_n8757_;
  assign new_n8764_ = new_n8295_ & new_n8729_;
  assign new_n5285_ = ~new_n8764_;
  assign new_n8769_ = new_n8794_ & new_n7536_;
  assign new_n5286_ = ~new_n8769_;
  assign new_n8771_ = new_n6091_ & new_n5801_;
  assign new_n5287_ = ~new_n8771_;
  assign new_n8782_ = new_n7998_ & new_n9269_;
  assign new_n7305_ = ~new_n9560_;
  assign new_n5288_ = ~new_n8782_;
  assign new_n8784_ = new_n8433_ & new_n8805_;
  assign new_n5289_ = ~new_n8784_;
  assign new_n8791_ = new_n8295_ & new_n8750_;
  assign new_n5290_ = ~new_n8791_;
  assign new_n8803_ = new_n8800_ & new_n7419_;
  assign new_n5291_ = ~new_n8803_;
  assign new_n8810_ = new_n8015_ & new_n9269_;
  assign new_n5292_ = ~new_n8810_;
  assign new_n8812_ = new_n8433_ & new_n8841_;
  assign new_n7055_ = ~new_n10525_;
  assign new_n7306_ = ~new_n9902_;
  assign new_n5293_ = ~new_n8812_;
  assign new_n8818_ = new_n6094_ & new_n7542_;
  assign new_n5294_ = ~new_n8818_;
  assign new_n8827_ = new_n8295_ & new_n8774_;
  assign new_n5295_ = ~new_n8827_;
  assign new_n8832_ = new_n8862_ & new_n7532_;
  assign new_n5296_ = ~new_n8832_;
  assign new_n8847_ = new_n8032_ & new_n9269_;
  assign new_n5297_ = ~new_n8847_;
  assign new_n8849_ = new_n8433_ & new_n8869_;
  assign new_n10436_ = new_n7456_ & new_n8750_;
  assign new_n5298_ = ~new_n8849_;
  assign new_n8855_ = new_n7356_ & new_n7470_;
  assign new_n5299_ = ~new_n8855_;
  assign new_n8859_ = new_n8295_ & new_n8805_;
  assign new_n5300_ = ~new_n8859_;
  assign new_n8864_ = new_n8865_ & new_n7282_;
  assign new_n5301_ = ~new_n8864_;
  assign new_n8866_ = new_n7156_ & new_n5805_;
  assign new_n5302_ = ~new_n8866_;
  assign new_n8874_ = new_n8049_ & new_n9269_;
  assign new_n7307_ = ~new_n10436_;
  assign new_n5303_ = ~new_n8874_;
  assign new_n8876_ = new_n8433_ & new_n8927_;
  assign new_n5304_ = ~new_n8876_;
  assign new_n8882_ = new_n8295_ & new_n8841_;
  assign new_n5305_ = ~new_n8882_;
  assign new_n8887_ = new_n8916_ & new_n7437_;
  assign new_n5306_ = ~new_n8887_;
  assign new_n8893_ = new_n8894_ & new_n7123_;
  assign new_n5307_ = ~new_n8893_;
  assign new_n8904_ = new_n8066_ & new_n9269_;
  assign new_n10686_ = new_n7528_ & new_n9405_;
  assign new_n5308_ = ~new_n8904_;
  assign new_n8906_ = new_n8433_ & new_n8928_;
  assign new_n5309_ = ~new_n8906_;
  assign new_n8913_ = new_n8295_ & new_n8869_;
  assign new_n5310_ = ~new_n8913_;
  assign new_n8925_ = new_n7123_ & new_n7436_;
  assign new_n5311_ = ~new_n8925_;
  assign new_n8933_ = new_n8083_ & new_n9269_;
  assign new_n5312_ = ~new_n8933_;
  assign new_n8935_ = new_n8433_ & new_n8952_;
  assign new_n7308_ = ~new_n10686_;
  assign new_n5313_ = ~new_n8935_;
  assign new_n8944_ = new_n8295_ & new_n8927_;
  assign new_n5314_ = ~new_n8944_;
  assign new_n8949_ = new_n8117_ & new_n7445_;
  assign new_n5315_ = ~new_n8949_;
  assign new_n8950_ = new_n8891_ & new_n5809_;
  assign new_n5316_ = ~new_n8950_;
  assign new_n8957_ = new_n8100_ & new_n9269_;
  assign new_n5317_ = ~new_n8957_;
  assign new_n8959_ = new_n8433_ & new_n9024_;
  assign new_n10664_ = new_n7396_ & new_n9419_;
  assign new_n5318_ = ~new_n8959_;
  assign new_n8965_ = new_n6103_ & new_n7399_;
  assign new_n5319_ = ~new_n8965_;
  assign new_n8974_ = new_n8295_ & new_n8928_;
  assign new_n5320_ = ~new_n8974_;
  assign new_n8978_ = new_n8979_ & new_n8989_;
  assign new_n5321_ = ~new_n8978_;
  assign new_n8994_ = new_n8119_ & new_n9269_;
  assign new_n5322_ = ~new_n8994_;
  assign new_n8996_ = new_n8433_ & new_n9025_;
  assign new_n7309_ = ~new_n10664_;
  assign new_n5323_ = ~new_n8996_;
  assign new_n8999_ = new_n6106_ & new_n9001_;
  assign new_n5324_ = ~new_n8999_;
  assign new_n9004_ = new_n7415_ & new_n7366_;
  assign new_n5325_ = ~new_n9004_;
  assign new_n9008_ = new_n8295_ & new_n8952_;
  assign new_n5326_ = ~new_n9008_;
  assign new_n9013_ = new_n8152_ & new_n7535_;
  assign new_n5327_ = ~new_n9013_;
  assign new_n9022_ = new_n7124_ & new_n7433_;
  assign new_n8624_ = new_n7479_ & new_n10496_;
  assign new_n5328_ = ~new_n9022_;
  assign new_n9030_ = new_n8136_ & new_n9269_;
  assign new_n5329_ = ~new_n9030_;
  assign new_n9032_ = new_n8433_ & new_n9043_;
  assign new_n5330_ = ~new_n9032_;
  assign new_n9038_ = new_n8295_ & new_n9024_;
  assign new_n5331_ = ~new_n9038_;
  assign new_n9041_ = new_n8981_ & new_n5814_;
  assign new_n5332_ = ~new_n9041_;
  assign new_n9048_ = new_n8154_ & new_n9269_;
  assign new_n7310_ = ~new_n8624_;
  assign new_n5333_ = ~new_n9048_;
  assign new_n9050_ = new_n8433_ & new_n9075_;
  assign new_n5334_ = ~new_n9050_;
  assign new_n9065_ = new_n8295_ & new_n9025_;
  assign new_n5335_ = ~new_n9065_;
  assign new_n9070_ = new_n8187_ & new_n7534_;
  assign new_n5336_ = ~new_n9070_;
  assign new_n9072_ = new_n6110_ & new_n5817_;
  assign new_n5337_ = ~new_n9072_;
  assign new_n9083_ = new_n8171_ & new_n9269_;
  assign new_n7311_ = ~new_n8835_;
  assign new_n5338_ = ~new_n9083_;
  assign new_n9085_ = new_n8433_ & new_n9106_;
  assign new_n5339_ = ~new_n9085_;
  assign new_n9093_ = new_n8295_ & new_n9043_;
  assign new_n5340_ = ~new_n9093_;
  assign new_n9104_ = new_n9101_ & new_n7420_;
  assign new_n5341_ = ~new_n9104_;
  assign new_n9105_ = new_n7371_ & new_n7534_;
  assign new_n5342_ = ~new_n9105_;
  assign new_n9111_ = new_n8189_ & new_n9269_;
  assign new_n7056_ = ~new_n10703_;
  assign new_n7312_ = ~new_n9804_;
  assign new_n5343_ = ~new_n9111_;
  assign new_n9113_ = new_n8433_ & new_n9173_;
  assign new_n5344_ = ~new_n9113_;
  assign new_n9128_ = new_n8295_ & new_n9075_;
  assign new_n5345_ = ~new_n9128_;
  assign new_n9134_ = new_n7429_ & new_n7533_;
  assign new_n5346_ = ~new_n9134_;
  assign new_n9146_ = new_n8206_ & new_n9269_;
  assign new_n5347_ = ~new_n9146_;
  assign new_n9148_ = new_n8433_ & new_n9171_;
  assign new_n11461_ = new_n9352_ & new_n9351_;
  assign new_n5348_ = ~new_n9148_;
  assign new_n9151_ = new_n6115_ & new_n9153_;
  assign new_n5349_ = ~new_n9151_;
  assign new_n9158_ = new_n8295_ & new_n9106_;
  assign new_n5350_ = ~new_n9158_;
  assign new_n9169_ = new_n9166_ & new_n7421_;
  assign new_n5351_ = ~new_n9169_;
  assign new_n9178_ = new_n9172_ & new_n9269_;
  assign new_n5352_ = ~new_n9178_;
  assign new_n9180_ = new_n8433_ & new_n8262_;
  assign new_n7313_ = ~new_n11461_;
  assign new_n5353_ = ~new_n9180_;
  assign new_n9187_ = new_n8295_ & new_n9173_;
  assign new_n5354_ = ~new_n9187_;
  assign new_n9194_ = new_n9195_ & new_n8262_;
  assign new_n5355_ = ~new_n9194_;
  assign new_n9201_ = new_n8239_ & new_n9269_;
  assign new_n5356_ = ~new_n9201_;
  assign new_n9203_ = new_n8433_ & new_n9216_;
  assign new_n5357_ = ~new_n9203_;
  assign new_n9210_ = new_n8295_ & new_n9171_;
  assign new_n7314_ = ~new_n10134_;
  assign new_n5358_ = ~new_n9210_;
  assign new_n9214_ = new_n7126_ & new_n5824_;
  assign new_n5359_ = ~new_n9214_;
  assign new_n9221_ = new_n8257_ & new_n9269_;
  assign new_n5360_ = ~new_n9221_;
  assign new_n9223_ = new_n8433_ & new_n10442_;
  assign new_n5361_ = ~new_n9223_;
  assign new_n9230_ = new_n8295_ & new_n8262_;
  assign new_n5362_ = ~new_n9230_;
  assign new_n9236_ = new_n7549_ & new_n7394_;
  assign new_n7315_ = ~new_n10006_;
  assign new_n5363_ = ~new_n9236_;
  assign new_n9249_ = new_n8274_ & new_n9269_;
  assign new_n5364_ = ~new_n9249_;
  assign new_n9251_ = new_n8433_ & new_n10586_;
  assign new_n5365_ = ~new_n9251_;
  assign new_n9258_ = new_n8295_ & new_n9216_;
  assign new_n5366_ = ~new_n9258_;
  assign new_n9264_ = new_n8295_ & new_n10442_;
  assign new_n5367_ = ~new_n9264_;
  assign new_n9268_ = new_n7265_ & new_n7256_;
  assign new_n7316_ = ~new_n10034_;
  assign new_n5368_ = ~new_n9268_;
  assign new_n9273_ = new_n7701_ & new_n9278_;
  assign new_n5369_ = ~new_n9273_;
  assign new_n9277_ = new_n10135_ & new_n7547_;
  assign new_n5370_ = ~new_n9277_;
  assign new_n9310_ = new_n7553_ & new_n9312_;
  assign new_n5371_ = ~new_n9310_;
  assign new_n9326_ = new_n7553_ & new_n5835_;
  assign new_n5372_ = ~new_n9326_;
  assign new_n9334_ = new_n7553_ & new_n5837_;
  assign new_n7317_ = ~new_n10055_;
  assign new_n5373_ = ~new_n9334_;
  assign new_n9348_ = new_n7553_ & new_n5840_;
  assign new_n5374_ = ~new_n9348_;
  assign new_n9357_ = new_n7553_ & new_n5842_;
  assign new_n5375_ = ~new_n9357_;
  assign new_n9372_ = new_n7553_ & new_n5845_;
  assign new_n5376_ = ~new_n9372_;
  assign new_n9387_ = new_n7553_ & new_n5848_;
  assign new_n5377_ = ~new_n9387_;
  assign new_n9401_ = new_n7553_ & new_n5851_;
  assign new_n7318_ = ~new_n10064_;
  assign new_n5378_ = ~new_n9401_;
  assign new_n9415_ = new_n7553_ & new_n5854_;
  assign new_n5379_ = ~new_n9415_;
  assign new_n9430_ = new_n7553_ & new_n5857_;
  assign new_n5380_ = ~new_n9430_;
  assign new_n9445_ = new_n7553_ & new_n5860_;
  assign new_n5381_ = ~new_n9445_;
  assign new_n9460_ = new_n7553_ & new_n5863_;
  assign new_n5382_ = ~new_n9460_;
  assign new_n9475_ = new_n7553_ & new_n5866_;
  assign new_n7319_ = ~new_n10043_;
  assign new_n5383_ = ~new_n9475_;
  assign new_n9490_ = new_n7553_ & new_n5869_;
  assign new_n5384_ = ~new_n9490_;
  assign new_n9504_ = new_n7553_ & new_n5872_;
  assign new_n5385_ = ~new_n9504_;
  assign new_n9513_ = new_n7553_ & new_n5874_;
  assign new_n5386_ = ~new_n9513_;
  assign new_n9528_ = new_n7553_ & new_n5877_;
  assign new_n5387_ = ~new_n9528_;
  assign new_n9546_ = new_n9547_ & new_n9106_;
  assign new_n7320_ = ~new_n10096_;
  assign new_n5388_ = ~new_n9546_;
  assign new_n9550_ = new_n8176_ & new_n7555_;
  assign new_n5389_ = ~new_n9550_;
  assign new_n9557_ = new_n9558_ & new_n5880_;
  assign new_n5390_ = ~new_n9557_;
  assign new_n9572_ = REG3_REG_27_ & n1332;
  assign new_n5391_ = ~new_n9572_;
  assign new_n9574_ = new_n9547_ & new_n8553_;
  assign new_n5392_ = ~new_n9574_;
  assign new_n9576_ = new_n7833_ & new_n7555_;
  assign new_n7608_ = new_n7729_ & new_n7120_;
  assign new_n7321_ = ~new_n10186_;
  assign new_n5393_ = ~new_n9576_;
  assign new_n9588_ = new_n9547_ & new_n8927_;
  assign new_n5394_ = ~new_n9588_;
  assign new_n9590_ = new_n7294_ & new_n7555_;
  assign new_n5395_ = ~new_n9590_;
  assign new_n9601_ = REG3_REG_23_ & n1332;
  assign new_n5396_ = ~new_n9601_;
  assign new_n9603_ = new_n9547_ & new_n8637_;
  assign new_n5397_ = ~new_n9603_;
  assign new_n9605_ = new_n7901_ & new_n7555_;
  assign new_n7322_ = ~new_n10196_;
  assign new_n5398_ = ~new_n9605_;
  assign new_n9618_ = new_n9547_ & new_n9025_;
  assign new_n5399_ = ~new_n9618_;
  assign new_n9620_ = new_n8124_ & new_n7555_;
  assign new_n5400_ = ~new_n9620_;
  assign new_n9630_ = new_n9548_ & new_n9171_;
  assign new_n5401_ = ~new_n9630_;
  assign new_n9634_ = new_n9547_ & new_n9216_;
  assign new_n5402_ = ~new_n9634_;
  assign new_n9653_ = new_n9547_ & new_n8750_;
  assign new_n7323_ = ~new_n10209_;
  assign new_n5403_ = ~new_n9653_;
  assign new_n9655_ = new_n7969_ & new_n7555_;
  assign new_n5404_ = ~new_n9655_;
  assign new_n9666_ = REG3_REG_28_ & n1332;
  assign new_n5405_ = ~new_n9666_;
  assign new_n9668_ = new_n9547_ & new_n8483_;
  assign new_n5406_ = ~new_n9668_;
  assign new_n9670_ = new_n7816_ & new_n7555_;
  assign new_n5407_ = ~new_n9670_;
  assign new_n9679_ = new_n7808_ & new_n7557_;
  assign new_n7324_ = ~new_n10220_;
  assign new_n5408_ = ~new_n9679_;
  assign new_n9683_ = new_n9681_ & new_n7808_;
  assign new_n5409_ = ~new_n9683_;
  assign new_n9687_ = new_n9581_ & new_n9688_;
  assign new_n5410_ = ~new_n9687_;
  assign new_n9691_ = new_n7828_ & new_n7557_;
  assign new_n5411_ = ~new_n9691_;
  assign new_n9703_ = new_n9547_ & new_n9075_;
  assign new_n5412_ = ~new_n9703_;
  assign new_n9705_ = new_n8159_ & new_n7555_;
  assign new_n7325_ = ~new_n10229_;
  assign new_n5413_ = ~new_n9705_;
  assign new_n9716_ = new_n9547_ & new_n10586_;
  assign new_n5414_ = ~new_n9716_;
  assign new_n9718_ = new_n8274_ & new_n7556_;
  assign new_n5415_ = ~new_n9718_;
  assign new_n9730_ = REG3_REG_21_ & n1332;
  assign new_n5416_ = ~new_n9730_;
  assign new_n9732_ = new_n9547_ & new_n8728_;
  assign new_n5417_ = ~new_n9732_;
  assign new_n9734_ = new_n7935_ & new_n7555_;
  assign new_n7326_ = ~new_n10242_;
  assign new_n5418_ = ~new_n9734_;
  assign new_n9739_ = new_n9740_ & new_n7202_;
  assign new_n5419_ = ~new_n9739_;
  assign new_n9754_ = new_n9547_ & new_n8952_;
  assign new_n5420_ = ~new_n9754_;
  assign new_n9756_ = new_n8088_ & new_n7555_;
  assign new_n5421_ = ~new_n9756_;
  assign new_n9766_ = REG3_REG_25_ & n1332;
  assign new_n5422_ = ~new_n9766_;
  assign new_n9768_ = new_n9547_ & new_n8521_;
  assign new_n7327_ = ~new_n10165_;
  assign new_n5423_ = ~new_n9768_;
  assign new_n9770_ = new_n7867_ & new_n7555_;
  assign new_n5424_ = ~new_n9770_;
  assign new_n9782_ = new_n9547_ & new_n8841_;
  assign new_n5425_ = ~new_n9782_;
  assign new_n9784_ = new_n8020_ & new_n7555_;
  assign new_n5426_ = ~new_n9784_;
  assign new_n9796_ = new_n9547_ & new_n9171_;
  assign new_n5427_ = ~new_n9796_;
  assign new_n9798_ = new_n8211_ & new_n7555_;
  assign new_n7328_ = ~new_n10151_;
  assign new_n5428_ = ~new_n9798_;
  assign new_n9809_ = new_n9547_ & new_n8805_;
  assign new_n5429_ = ~new_n9809_;
  assign new_n9811_ = new_n8003_ & new_n7555_;
  assign new_n5430_ = ~new_n9811_;
  assign new_n9816_ = new_n9817_ & new_n7203_;
  assign new_n5431_ = ~new_n9816_;
  assign new_n9827_ = REG3_REG_24_ & n1332;
  assign new_n5432_ = ~new_n9827_;
  assign new_n9829_ = new_n9547_ & new_n8596_;
  assign new_n7329_ = ~new_n10157_;
  assign new_n5433_ = ~new_n9829_;
  assign new_n9831_ = new_n7884_ & new_n7555_;
  assign new_n5434_ = ~new_n9831_;
  assign new_n9844_ = new_n9547_ & new_n8262_;
  assign new_n5435_ = ~new_n9844_;
  assign new_n9846_ = new_n9172_ & new_n7556_;
  assign new_n5436_ = ~new_n9846_;
  assign new_n9859_ = new_n9547_ & new_n9043_;
  assign new_n5437_ = ~new_n9859_;
  assign new_n9861_ = new_n8141_ & new_n7555_;
  assign new_n7330_ = ~new_n8671_;
  assign new_n5438_ = ~new_n9861_;
  assign new_n9872_ = new_n9554_ & new_n9873_;
  assign new_n5439_ = ~new_n9872_;
  assign new_n9875_ = REG3_REG_0_ & new_n9726_;
  assign new_n5440_ = ~new_n9875_;
  assign new_n9879_ = REG3_REG_20_ & n1332;
  assign new_n5441_ = ~new_n9879_;
  assign new_n9881_ = new_n9547_ & new_n8729_;
  assign new_n5442_ = ~new_n9881_;
  assign new_n9883_ = new_n7952_ & new_n7555_;
  assign new_n7057_ = ~new_n7608_;
  assign new_n7331_ = ~new_n7708_;
  assign new_n5443_ = ~new_n9883_;
  assign new_n9892_ = new_n9547_ & new_n8928_;
  assign new_n5444_ = ~new_n9892_;
  assign new_n9894_ = new_n8071_ & new_n7555_;
  assign new_n5445_ = ~new_n9894_;
  assign new_n9901_ = new_n7306_ & new_n7274_;
  assign new_n5446_ = ~new_n9901_;
  assign new_n9910_ = new_n7158_ & new_n7441_;
  assign new_n5447_ = ~new_n9910_;
  assign new_n9916_ = REG3_REG_22_ & n1332;
  assign new_n7332_ = ~new_n7706_;
  assign new_n5448_ = ~new_n9916_;
  assign new_n9918_ = new_n9547_ & new_n8674_;
  assign new_n5449_ = ~new_n9918_;
  assign new_n9920_ = new_n7293_ & new_n7555_;
  assign new_n5450_ = ~new_n9920_;
  assign new_n9933_ = new_n9547_ & new_n9024_;
  assign new_n5451_ = ~new_n9933_;
  assign new_n9935_ = new_n8105_ & new_n7555_;
  assign new_n5452_ = ~new_n9935_;
  assign new_n9938_ = new_n9939_ & new_n9940_;
  assign new_n7333_ = ~new_n8800_;
  assign new_n5453_ = ~new_n9938_;
  assign new_n9947_ = new_n7291_ & new_n7037_;
  assign new_n5454_ = ~new_n9947_;
  assign new_n9952_ = new_n9547_ & new_n10442_;
  assign new_n5455_ = ~new_n9952_;
  assign new_n9954_ = new_n8257_ & new_n7556_;
  assign new_n5456_ = ~new_n9954_;
  assign new_n9963_ = new_n9547_ & new_n8774_;
  assign new_n5457_ = ~new_n9963_;
  assign new_n9965_ = new_n7986_ & new_n7555_;
  assign new_n8800_ = new_n8833_ & new_n8834_;
  assign new_n5458_ = ~new_n9965_;
  assign new_n9978_ = new_n9547_ & new_n9173_;
  assign new_n5459_ = ~new_n9978_;
  assign new_n9980_ = new_n8194_ & new_n7555_;
  assign new_n5460_ = ~new_n9980_;
  assign new_n9985_ = new_n7312_ & new_n7038_;
  assign new_n5461_ = ~new_n9985_;
  assign new_n9990_ = REG3_REG_26_ & n1332;
  assign new_n5462_ = ~new_n9990_;
  assign new_n9992_ = new_n9547_ & new_n8552_;
  assign new_n7334_ = ~new_n9101_;
  assign new_n5463_ = ~new_n9992_;
  assign new_n9994_ = new_n7850_ & new_n7555_;
  assign new_n5464_ = ~new_n9994_;
  assign new_n10009_ = new_n9681_ & new_n7862_;
  assign new_n5465_ = ~new_n10009_;
  assign new_n10011_ = new_n7862_ & new_n7557_;
  assign new_n5466_ = ~new_n10011_;
  assign new_n10013_ = new_n9835_ & new_n10014_;
  assign new_n5467_ = ~new_n10013_;
  assign new_n10017_ = new_n7879_ & new_n7557_;
  assign new_n9101_ = new_n9135_ & new_n9136_;
  assign new_n5468_ = ~new_n10017_;
  assign new_n10019_ = new_n9681_ & new_n7879_;
  assign new_n5469_ = ~new_n10019_;
  assign new_n10021_ = new_n9609_ & new_n10022_;
  assign new_n5470_ = ~new_n10021_;
  assign new_n10025_ = new_n7896_ & new_n7557_;
  assign new_n5471_ = ~new_n10025_;
  assign new_n10027_ = new_n9681_ & new_n7896_;
  assign new_n5472_ = ~new_n10027_;
  assign new_n10029_ = new_n9926_ & new_n10030_;
  assign new_n7335_ = ~new_n8667_;
  assign new_n5473_ = ~new_n10029_;
  assign new_n10037_ = new_n9681_ & new_n7930_;
  assign new_n5474_ = ~new_n10037_;
  assign new_n10039_ = new_n7930_ & new_n7557_;
  assign new_n5475_ = ~new_n10039_;
  assign new_n10045_ = new_n9662_ & new_n5881_;
  assign new_n5476_ = ~new_n10045_;
  assign new_n10058_ = new_n9681_ & new_n7998_;
  assign new_n5477_ = ~new_n10058_;
  assign new_n10060_ = new_n7998_ & new_n7557_;
  assign new_n7336_ = ~new_n8891_;
  assign new_n5478_ = ~new_n10060_;
  assign new_n10066_ = new_n6144_ & new_n7221_;
  assign new_n5479_ = ~new_n10066_;
  assign new_n10073_ = new_n9681_ & new_n8015_;
  assign new_n5480_ = ~new_n10073_;
  assign new_n10075_ = new_n8015_ & new_n7557_;
  assign new_n5481_ = ~new_n10075_;
  assign new_n10078_ = new_n7981_ & new_n7557_;
  assign new_n5482_ = ~new_n10078_;
  assign new_n10080_ = new_n9681_ & new_n7981_;
  assign new_n7337_ = ~new_n8981_;
  assign new_n5483_ = ~new_n10080_;
  assign new_n10083_ = new_n7964_ & new_n7557_;
  assign new_n5484_ = ~new_n10083_;
  assign new_n10086_ = new_n9681_ & new_n7947_;
  assign new_n5485_ = ~new_n10086_;
  assign new_n10088_ = new_n7947_ & new_n7557_;
  assign new_n5486_ = ~new_n10088_;
  assign new_n10090_ = new_n9681_ & new_n7913_;
  assign new_n5487_ = ~new_n10090_;
  assign new_n10093_ = new_n7913_ & new_n7557_;
  assign new_n7338_ = ~new_n10740_;
  assign new_n5488_ = ~new_n10093_;
  assign new_n10099_ = new_n9681_ & new_n7845_;
  assign new_n5489_ = ~new_n10099_;
  assign new_n10101_ = new_n7845_ & new_n7557_;
  assign new_n5490_ = ~new_n10101_;
  assign new_n10106_ = new_n9547_ & new_n8869_;
  assign new_n5491_ = ~new_n10106_;
  assign new_n10111_ = new_n8037_ & new_n7555_;
  assign new_n5492_ = ~new_n10111_;
  assign new_n10113_ = new_n10114_ & new_n10703_;
  assign new_n8892_ = new_n7246_ & new_n7437_;
  assign new_n10740_ = new_n10758_ & REG3_REG_26_;
  assign new_n5493_ = ~new_n10113_;
  assign new_n10120_ = new_n7187_ & new_n10122_;
  assign new_n5494_ = ~new_n10120_;
  assign new_n10129_ = new_n8413_ & new_n7545_;
  assign new_n5495_ = ~new_n10129_;
  assign new_n10142_ = new_n8032_ & new_n7557_;
  assign new_n5496_ = ~new_n10142_;
  assign new_n10144_ = new_n9681_ & new_n8032_;
  assign new_n5497_ = ~new_n10144_;
  assign new_n10146_ = new_n6147_ & new_n7222_;
  assign new_n10761_ = new_n10779_ & REG3_REG_24_;
  assign new_n5498_ = ~new_n10146_;
  assign new_n10160_ = new_n9909_ & new_n5883_;
  assign new_n5499_ = ~new_n10160_;
  assign new_n10167_ = new_n9867_ & new_n5885_;
  assign new_n5500_ = ~new_n10167_;
  assign new_n10179_ = new_n9853_ & new_n5886_;
  assign new_n5501_ = ~new_n10179_;
  assign new_n10189_ = new_n9681_ & new_n8239_;
  assign new_n5502_ = ~new_n10189_;
  assign new_n10191_ = new_n8239_ & new_n7557_;
  assign new_n7339_ = ~new_n10761_;
  assign new_n5503_ = ~new_n10191_;
  assign new_n10193_ = new_n7228_ & new_n7134_;
  assign new_n5504_ = ~new_n10193_;
  assign new_n10198_ = new_n10199_ & new_n7569_;
  assign new_n5505_ = ~new_n10198_;
  assign new_n10204_ = new_n9681_ & new_n8274_;
  assign new_n5506_ = ~new_n10204_;
  assign new_n10206_ = new_n8274_ & new_n7557_;
  assign new_n5507_ = ~new_n10206_;
  assign new_n10212_ = new_n9681_ & new_n8257_;
  assign new_n10843_ = new_n10861_ & new_n7440_;
  assign new_n5508_ = ~new_n10212_;
  assign new_n10214_ = new_n8257_ & new_n7557_;
  assign new_n5509_ = ~new_n10214_;
  assign new_n10217_ = new_n9172_ & new_n7557_;
  assign new_n5510_ = ~new_n10217_;
  assign new_n10223_ = new_n8206_ & new_n7557_;
  assign new_n5511_ = ~new_n10223_;
  assign new_n10225_ = new_n9681_ & new_n8206_;
  assign new_n5512_ = ~new_n10225_;
  assign new_n10232_ = new_n9681_ & new_n8189_;
  assign new_n7340_ = ~new_n10843_;
  assign new_n5513_ = ~new_n10232_;
  assign new_n10234_ = new_n8189_ & new_n7557_;
  assign new_n5514_ = ~new_n10234_;
  assign new_n10237_ = new_n9681_ & new_n8171_;
  assign new_n5515_ = ~new_n10237_;
  assign new_n10239_ = new_n8171_ & new_n7557_;
  assign new_n5516_ = ~new_n10239_;
  assign new_n10245_ = new_n9681_ & new_n8154_;
  assign new_n5517_ = ~new_n10245_;
  assign new_n10247_ = new_n8154_ & new_n7557_;
  assign new_n10905_ = new_n10923_ & REG3_REG_9_;
  assign new_n5518_ = ~new_n10247_;
  assign new_n10250_ = new_n8136_ & new_n7557_;
  assign new_n5519_ = ~new_n10250_;
  assign new_n10252_ = new_n9681_ & new_n8136_;
  assign new_n5520_ = ~new_n10252_;
  assign new_n10255_ = new_n9681_ & new_n8119_;
  assign new_n5521_ = ~new_n10255_;
  assign new_n10257_ = new_n8119_ & new_n7557_;
  assign new_n5522_ = ~new_n10257_;
  assign new_n10259_ = new_n9681_ & new_n8100_;
  assign new_n7341_ = ~new_n10905_;
  assign new_n5523_ = ~new_n10259_;
  assign new_n10262_ = new_n8100_ & new_n7557_;
  assign new_n5524_ = ~new_n10262_;
  assign new_n10265_ = new_n9681_ & new_n8066_;
  assign new_n5525_ = ~new_n10265_;
  assign new_n10267_ = new_n8066_ & new_n7557_;
  assign new_n5526_ = ~new_n10267_;
  assign new_n5527_ = ~new_n10155_;
  assign new_n10270_ = new_n8083_ & new_n7557_;
  assign new_n5528_ = ~new_n10270_;
  assign new_n10926_ = new_n10944_ & REG3_REG_8_;
  assign new_n10273_ = new_n8049_ & new_n7557_;
  assign new_n5529_ = ~new_n10273_;
  assign new_n10275_ = new_n9681_ & new_n8049_;
  assign new_n5530_ = ~new_n10275_;
  assign new_n10276_ = new_n10277_ & new_n7230_;
  assign new_n5531_ = ~new_n10276_;
  assign new_n10280_ = new_n7196_ & new_n10281_;
  assign new_n5532_ = ~new_n10280_;
  assign new_n10286_ = new_n9300_ & new_n5888_;
  assign new_n5533_ = ~new_n10286_;
  assign new_n7342_ = ~new_n10926_;
  assign new_n10301_ = new_n9300_ & new_n5892_;
  assign new_n5534_ = ~new_n10301_;
  assign new_n10335_ = new_n6152_ & new_n7469_;
  assign new_n5535_ = ~new_n10335_;
  assign new_n10339_ = new_n10340_ & new_n5898_;
  assign new_n5536_ = ~new_n10339_;
  assign new_n10373_ = new_n10374_ & new_n10375_;
  assign new_n5537_ = ~new_n10373_;
  assign new_n10387_ = new_n10388_ & new_n10389_;
  assign new_n5538_ = ~new_n10387_;
  assign new_n7343_ = ~new_n10966_;
  assign new_n10408_ = new_n10409_ & new_n10405_;
  assign new_n5539_ = ~new_n10408_;
  assign new_n10425_ = new_n6294_ | new_n6703_;
  assign new_n5540_ = ~new_n10425_;
  assign new_n10429_ = new_n6292_ | new_n6704_;
  assign new_n5541_ = ~new_n10429_;
  assign new_n10438_ = new_n6295_ | new_n7214_;
  assign new_n5542_ = ~new_n10438_;
  assign new_n10449_ = new_n6297_ | new_n6708_;
  assign new_n5543_ = ~new_n10449_;
  assign new_n7058_ = ~new_n8892_;
  assign new_n10966_ = REG3_REG_4_ & REG3_REG_3_;
  assign new_n10457_ = new_n6300_ | new_n6709_;
  assign new_n5544_ = ~new_n10457_;
  assign new_n10469_ = new_n10138_ & new_n10470_;
  assign new_n5545_ = ~new_n10469_;
  assign new_n10474_ = new_n10478_ & new_n5914_;
  assign new_n5546_ = ~new_n10474_;
  assign new_n10477_ = new_n7413_ & new_n7514_;
  assign new_n5547_ = ~new_n10477_;
  assign new_n10481_ = new_n10445_ & new_n7110_;
  assign new_n5548_ = ~new_n10481_;
  assign new_n7344_ = ~new_n8444_;
  assign new_n10490_ = new_n7522_ & new_n7205_;
  assign new_n5549_ = ~new_n10490_;
  assign new_n10492_ = new_n6160_ & new_n7482_;
  assign new_n5550_ = ~new_n10492_;
  assign new_n10494_ = new_n8629_ & new_n7530_;
  assign new_n5551_ = ~new_n10494_;
  assign new_n10499_ = new_n7406_ & new_n7225_;
  assign new_n5552_ = ~new_n10499_;
  assign new_n10500_ = new_n7223_ & new_n7409_;
  assign new_n5553_ = ~new_n10500_;
  assign new_n7345_ = ~new_n9775_;
  assign new_n10502_ = new_n6161_ & new_n7452_;
  assign new_n5554_ = ~new_n10502_;
  assign new_n10505_ = new_n8854_ & new_n7541_;
  assign new_n5555_ = ~new_n10505_;
  assign new_n10508_ = new_n8910_ & new_n7302_;
  assign new_n5556_ = ~new_n10508_;
  assign new_n10513_ = new_n9090_ & new_n10390_;
  assign new_n5557_ = ~new_n10513_;
  assign new_n10524_ = new_n7549_ & new_n7506_;
  assign new_n5558_ = ~new_n10524_;
  assign new_n7346_ = ~new_n9646_;
  assign new_n10526_ = new_n10384_ & new_n10383_;
  assign new_n5559_ = ~new_n10526_;
  assign new_n10528_ = new_n7480_ & new_n7521_;
  assign new_n5560_ = ~new_n10528_;
  assign new_n10530_ = new_n10324_ & new_n7045_;
  assign new_n5561_ = ~new_n10530_;
  assign new_n10535_ = new_n6303_ | new_n6713_;
  assign new_n5562_ = ~new_n10535_;
  assign new_n10543_ = new_n10544_ & new_n5919_;
  assign new_n5563_ = ~new_n10543_;
  assign new_n8685_ = new_n7526_ & new_n7546_;
  assign new_n10550_ = new_n6163_ & new_n7476_;
  assign new_n5564_ = ~new_n10550_;
  assign new_n10552_ = new_n10553_ & new_n7389_;
  assign new_n5565_ = ~new_n10552_;
  assign new_n10559_ = new_n7472_ & new_n5923_;
  assign new_n5566_ = ~new_n10559_;
  assign new_n10567_ = new_n10415_ & new_n7486_;
  assign new_n5567_ = ~new_n10567_;
  assign new_n10570_ = new_n7541_ & new_n5924_;
  assign new_n5568_ = ~new_n10570_;
  assign new_n7347_ = ~new_n8685_;
  assign new_n10573_ = new_n7054_ & new_n7515_;
  assign new_n5569_ = ~new_n10573_;
  assign new_n10574_ = new_n10464_ & new_n7529_;
  assign new_n5570_ = ~new_n10574_;
  assign new_n10585_ = new_n7550_ & new_n7506_;
  assign new_n5571_ = ~new_n10585_;
  assign new_n10623_ = new_n7303_ & new_n5928_;
  assign new_n5572_ = ~new_n10623_;
  assign new_n10627_ = new_n6167_ & new_n7388_;
  assign new_n5573_ = ~new_n10627_;
  assign new_n7348_ = ~new_n11248_;
  assign new_n10629_ = new_n6168_ & new_n7392_;
  assign new_n5574_ = ~new_n10629_;
  assign new_n10631_ = new_n8472_ & new_n7524_;
  assign new_n5575_ = ~new_n10631_;
  assign new_n10642_ = new_n10416_ & new_n7546_;
  assign new_n5576_ = ~new_n10642_;
  assign new_n10654_ = new_n6309_ | new_n6718_;
  assign new_n5577_ = ~new_n10654_;
  assign new_n10708_ = REG1_REG_31_ & new_n10709_;
  assign new_n5578_ = ~new_n10708_;
  assign new_n7349_ = ~new_n11090_;
  assign new_n10718_ = REG1_REG_30_ & new_n10709_;
  assign new_n5579_ = ~new_n10718_;
  assign new_n10726_ = REG2_REG_29_ & new_n7563_;
  assign new_n5580_ = ~new_n10726_;
  assign new_n10728_ = new_n10729_ & new_n7797_;
  assign new_n5581_ = ~new_n10728_;
  assign new_n10736_ = REG2_REG_28_ & new_n7563_;
  assign new_n5582_ = ~new_n10736_;
  assign new_n10738_ = new_n10729_ & new_n7816_;
  assign new_n5583_ = ~new_n10738_;
  assign new_n7350_ = ~new_n7738_;
  assign new_n10746_ = REG2_REG_27_ & new_n7563_;
  assign new_n5584_ = ~new_n10746_;
  assign new_n10748_ = new_n10729_ & new_n7833_;
  assign new_n5585_ = ~new_n10748_;
  assign new_n10754_ = REG2_REG_26_ & new_n7563_;
  assign new_n5586_ = ~new_n10754_;
  assign new_n10756_ = new_n7850_ & new_n10729_;
  assign new_n5587_ = ~new_n10756_;
  assign new_n10760_ = REG3_REG_25_ & new_n10761_;
  assign new_n5588_ = ~new_n10760_;
  assign new_n7783_ = new_n8414_ & new_n8449_;
  assign new_n10767_ = REG2_REG_25_ & new_n7563_;
  assign new_n5589_ = ~new_n10767_;
  assign new_n10769_ = new_n10729_ & new_n7867_;
  assign new_n5590_ = ~new_n10769_;
  assign new_n10775_ = REG2_REG_24_ & new_n7563_;
  assign new_n5591_ = ~new_n10775_;
  assign new_n10777_ = new_n7884_ & new_n10729_;
  assign new_n5592_ = ~new_n10777_;
  assign new_n10782_ = REG3_REG_23_ & new_n7439_;
  assign new_n5593_ = ~new_n10782_;
  assign new_n7059_ = ~new_n8398_;
  assign new_n7351_ = ~new_n7783_;
  assign new_n10788_ = REG2_REG_23_ & new_n7563_;
  assign new_n5594_ = ~new_n10788_;
  assign new_n10790_ = new_n10729_ & new_n7901_;
  assign new_n5595_ = ~new_n10790_;
  assign new_n10796_ = REG2_REG_22_ & new_n7563_;
  assign new_n5596_ = ~new_n10796_;
  assign new_n10798_ = new_n7293_ & new_n10729_;
  assign new_n5597_ = ~new_n10798_;
  assign new_n10807_ = REG2_REG_21_ & new_n7563_;
  assign new_n5598_ = ~new_n10807_;
  assign new_n7352_ = ~new_n8439_;
  assign new_n10809_ = new_n10729_ & new_n7935_;
  assign new_n5599_ = ~new_n10809_;
  assign new_n10816_ = REG2_REG_20_ & new_n7563_;
  assign new_n5600_ = ~new_n10816_;
  assign new_n10818_ = new_n7952_ & new_n10729_;
  assign new_n5601_ = ~new_n10818_;
  assign new_n5602_ = ~new_n10820_;
  assign new_n10828_ = new_n7563_ & REG2_REG_19_;
  assign new_n5603_ = ~new_n10828_;
  assign new_n10830_ = new_n10729_ & new_n7969_;
  assign new_n8439_ = new_n10420_ & new_n7392_;
  assign new_n5604_ = ~new_n10830_;
  assign new_n10836_ = new_n7563_ & REG2_REG_18_;
  assign new_n5605_ = ~new_n10836_;
  assign new_n10838_ = new_n7986_ & new_n10729_;
  assign new_n5606_ = ~new_n10838_;
  assign new_n10842_ = new_n10843_ & REG3_REG_17_;
  assign new_n5607_ = ~new_n10842_;
  assign new_n10849_ = new_n7563_ & REG2_REG_17_;
  assign new_n5608_ = ~new_n10849_;
  assign new_n10851_ = new_n10729_ & new_n8003_;
  assign new_n7353_ = ~new_n7626_;
  assign new_n5609_ = ~new_n10851_;
  assign new_n10857_ = new_n7563_ & REG2_REG_16_;
  assign new_n5610_ = ~new_n10857_;
  assign new_n10859_ = new_n8020_ & new_n10729_;
  assign new_n5611_ = ~new_n10859_;
  assign new_n10864_ = new_n7440_ & REG3_REG_15_;
  assign new_n5612_ = ~new_n10864_;
  assign new_n10870_ = new_n7563_ & REG2_REG_15_;
  assign new_n5613_ = ~new_n10870_;
  assign new_n10872_ = new_n10729_ & new_n8037_;
  assign new_n7354_ = ~new_n7587_;
  assign new_n5614_ = ~new_n10872_;
  assign new_n10878_ = new_n7563_ & REG2_REG_14_;
  assign new_n5615_ = ~new_n10878_;
  assign new_n10880_ = new_n7294_ & new_n10729_;
  assign new_n5616_ = ~new_n10880_;
  assign new_n10890_ = new_n7563_ & REG2_REG_13_;
  assign new_n5617_ = ~new_n10890_;
  assign new_n10892_ = new_n10729_ & new_n8071_;
  assign new_n5618_ = ~new_n10892_;
  assign new_n10898_ = REG2_REG_12_ & new_n7563_;
  assign new_n7355_ = ~new_n10822_;
  assign new_n5619_ = ~new_n10898_;
  assign new_n10900_ = new_n8088_ & new_n10729_;
  assign new_n5620_ = ~new_n10900_;
  assign new_n10904_ = REG3_REG_11_ & new_n10905_;
  assign new_n5621_ = ~new_n10904_;
  assign new_n10911_ = REG2_REG_11_ & new_n7563_;
  assign new_n5622_ = ~new_n10911_;
  assign new_n10913_ = new_n10729_ & new_n8105_;
  assign new_n5623_ = ~new_n10913_;
  assign new_n10919_ = REG2_REG_10_ & new_n7563_;
  assign new_n10822_ = new_n10840_ & new_n10843_;
  assign new_n5624_ = ~new_n10919_;
  assign new_n10921_ = new_n8124_ & new_n10729_;
  assign new_n5625_ = ~new_n10921_;
  assign new_n10925_ = REG3_REG_9_ & new_n10926_;
  assign new_n5626_ = ~new_n10925_;
  assign new_n10932_ = REG2_REG_9_ & new_n7563_;
  assign new_n5627_ = ~new_n10932_;
  assign new_n10934_ = new_n10729_ & new_n8141_;
  assign new_n5628_ = ~new_n10934_;
  assign new_n10940_ = REG2_REG_8_ & new_n7563_;
  assign new_n7356_ = ~new_n8856_;
  assign new_n5629_ = ~new_n10940_;
  assign new_n10942_ = new_n8159_ & new_n10729_;
  assign new_n5630_ = ~new_n10942_;
  assign new_n10947_ = REG3_REG_7_ & new_n10945_;
  assign new_n5631_ = ~new_n10947_;
  assign new_n10953_ = REG2_REG_7_ & new_n7563_;
  assign new_n5632_ = ~new_n10953_;
  assign new_n10955_ = new_n10729_ & new_n8176_;
  assign new_n5633_ = ~new_n10955_;
  assign new_n10962_ = REG2_REG_6_ & new_n7563_;
  assign new_n7357_ = ~new_n7610_;
  assign new_n5634_ = ~new_n10962_;
  assign new_n10964_ = new_n10729_ & new_n8194_;
  assign new_n5635_ = ~new_n10964_;
  assign new_n10972_ = REG2_REG_5_ & new_n7563_;
  assign new_n5636_ = ~new_n10972_;
  assign new_n10974_ = new_n10729_ & new_n8211_;
  assign new_n5637_ = ~new_n10974_;
  assign new_n10980_ = REG2_REG_4_ & new_n7563_;
  assign new_n5638_ = ~new_n10980_;
  assign new_n10982_ = new_n8222_ & new_n10729_;
  assign new_n7358_ = ~new_n8598_;
  assign new_n5639_ = ~new_n10982_;
  assign new_n10989_ = REG2_REG_3_ & new_n7563_;
  assign new_n5640_ = ~new_n10989_;
  assign new_n10991_ = REG0_REG_3_ & new_n7562_;
  assign new_n5641_ = ~new_n10991_;
  assign new_n10997_ = REG2_REG_2_ & new_n7563_;
  assign new_n5642_ = ~new_n10997_;
  assign new_n10999_ = REG0_REG_2_ & new_n7562_;
  assign new_n5643_ = ~new_n10999_;
  assign new_n11005_ = REG2_REG_1_ & new_n7563_;
  assign new_n11269_ = new_n11362_ & REG1_REG_10_;
  assign new_n7359_ = ~new_n9837_;
  assign new_n5644_ = ~new_n11005_;
  assign new_n11007_ = REG0_REG_1_ & new_n7562_;
  assign new_n5645_ = ~new_n11007_;
  assign new_n11013_ = ADDR_REG_0_ & new_n11294_;
  assign new_n5646_ = ~new_n11013_;
  assign new_n11027_ = ADDR_REG_1_ & new_n11294_;
  assign new_n5647_ = ~new_n11027_;
  assign new_n11043_ = REG3_REG_2_ & n1332;
  assign new_n5648_ = ~new_n11043_;
  assign new_n11045_ = new_n7446_ & new_n5965_;
  assign new_n7360_ = ~new_n9611_;
  assign new_n5649_ = ~new_n11045_;
  assign new_n11063_ = ADDR_REG_3_ & new_n11294_;
  assign new_n5650_ = ~new_n11063_;
  assign new_n11065_ = new_n7262_ & new_n5969_;
  assign new_n5651_ = ~new_n11065_;
  assign new_n11085_ = new_n10593_ & new_n5971_;
  assign new_n5652_ = ~new_n11085_;
  assign new_n11097_ = new_n7586_ & new_n11098_;
  assign new_n5653_ = ~new_n11097_;
  assign new_n11101_ = new_n6208_ & new_n7206_;
  assign new_n7361_ = ~new_n8485_;
  assign new_n5654_ = ~new_n11101_;
  assign new_n11111_ = IR_REG_0_ & new_n9540_;
  assign new_n5655_ = ~new_n11111_;
  assign new_n11121_ = REG1_REG_0_ & new_n9540_;
  assign new_n5656_ = ~new_n11121_;
  assign new_n11125_ = new_n6209_ & new_n9272_;
  assign new_n5657_ = ~new_n11125_;
  assign new_n11131_ = new_n10635_ & new_n9530_;
  assign new_n5658_ = ~new_n11131_;
  assign new_n11135_ = new_n7563_ & REG2_REG_0_;
  assign new_n7362_ = ~new_n8639_;
  assign new_n5659_ = ~new_n11135_;
  assign new_n11140_ = REG0_REG_0_ & new_n7562_;
  assign new_n5660_ = ~new_n11140_;
  assign new_n11142_ = IR_REG_29_ & new_n9536_;
  assign new_n5661_ = ~new_n11142_;
  assign new_n11156_ = ADDR_REG_5_ & new_n11294_;
  assign new_n5662_ = ~new_n11156_;
  assign new_n11158_ = new_n7261_ & new_n5973_;
  assign new_n5663_ = ~new_n11158_;
  assign new_n11176_ = ADDR_REG_6_ & new_n11294_;
  assign new_n7363_ = ~new_n9196_;
  assign new_n5664_ = ~new_n11176_;
  assign new_n11178_ = new_n7402_ & new_n5976_;
  assign new_n5665_ = ~new_n11178_;
  assign new_n11191_ = new_n7586_ & new_n11192_;
  assign new_n5666_ = ~new_n11191_;
  assign new_n11197_ = ADDR_REG_7_ & new_n11294_;
  assign new_n5667_ = ~new_n11197_;
  assign new_n11199_ = new_n7517_ & new_n5978_;
  assign new_n5668_ = ~new_n11199_;
  assign new_n11216_ = ADDR_REG_8_ & new_n11294_;
  assign new_n11033_ = REG2_REG_0_ & IR_REG_0_;
  assign new_n5669_ = ~new_n11216_;
  assign new_n11218_ = new_n10611_ & new_n5982_;
  assign new_n5670_ = ~new_n11218_;
  assign new_n11235_ = ADDR_REG_9_ & new_n11294_;
  assign new_n5671_ = ~new_n11235_;
  assign new_n11237_ = new_n7516_ & new_n5984_;
  assign new_n5672_ = ~new_n11237_;
  assign new_n11254_ = ADDR_REG_10_ & new_n11294_;
  assign new_n5673_ = ~new_n11254_;
  assign new_n11256_ = new_n10649_ & new_n5988_;
  assign new_n7364_ = ~new_n11033_;
  assign new_n5674_ = ~new_n11256_;
  assign new_n11273_ = ADDR_REG_11_ & new_n11294_;
  assign new_n5675_ = ~new_n11273_;
  assign new_n11275_ = new_n7460_ & new_n5990_;
  assign new_n5676_ = ~new_n11275_;
  assign new_n11293_ = ADDR_REG_12_ & new_n11294_;
  assign new_n5677_ = ~new_n11293_;
  assign new_n11296_ = new_n7739_ & new_n5994_;
  assign new_n5678_ = ~new_n11296_;
  assign new_n11309_ = new_n7586_ & new_n11310_;
  assign new_n7365_ = ~new_n8714_;
  assign new_n5679_ = ~new_n11309_;
  assign new_n11312_ = new_n11313_ & new_n11290_;
  assign new_n5680_ = ~new_n11312_;
  assign new_n11315_ = new_n11316_ & new_n11264_;
  assign new_n5681_ = ~new_n11315_;
  assign new_n11318_ = new_n11319_ & new_n11251_;
  assign new_n5682_ = ~new_n11318_;
  assign new_n11321_ = new_n11322_ & new_n11226_;
  assign new_n5683_ = ~new_n11321_;
  assign new_n11324_ = new_n11325_ & new_n11213_;
  assign new_n7366_ = ~new_n9006_;
  assign new_n5684_ = ~new_n11324_;
  assign new_n11327_ = new_n11328_ & new_n11188_;
  assign new_n5685_ = ~new_n11327_;
  assign new_n11330_ = new_n11331_ & new_n11167_;
  assign new_n5686_ = ~new_n11330_;
  assign new_n11333_ = new_n11334_ & new_n11094_;
  assign new_n5687_ = ~new_n11333_;
  assign new_n11336_ = new_n11337_ & new_n11074_;
  assign new_n5688_ = ~new_n11336_;
  assign new_n11339_ = new_n6222_ & new_n11050_;
  assign new_n7367_ = ~new_n8456_;
  assign new_n5689_ = ~new_n11339_;
  assign new_n11343_ = new_n11344_ & new_n11035_;
  assign new_n5690_ = ~new_n11343_;
  assign new_n11348_ = new_n6224_ & new_n11283_;
  assign new_n5691_ = ~new_n11348_;
  assign new_n11353_ = new_n10649_ & new_n7077_;
  assign new_n5692_ = ~new_n11353_;
  assign new_n11369_ = new_n10611_ & new_n7078_;
  assign new_n5693_ = ~new_n11369_;
  assign new_n11380_ = new_n7145_ & new_n11206_;
  assign new_n7026_ = ~new_n8127_;
  assign new_n7060_ = ~new_n11269_;
  assign new_n7368_ = ~new_n9582_;
  assign new_n5694_ = ~new_n11380_;
  assign new_n11383_ = new_n6227_ & new_n11194_;
  assign new_n5695_ = ~new_n11383_;
  assign new_n11387_ = new_n9536_ & new_n9494_;
  assign new_n5696_ = ~new_n11387_;
  assign new_n11389_ = new_n7261_ & new_n7079_;
  assign new_n5697_ = ~new_n11389_;
  assign new_n11395_ = IR_REG_5_ & new_n9536_;
  assign new_n5698_ = ~new_n11395_;
  assign new_n11405_ = new_n7262_ & new_n7080_;
  assign new_n7369_ = ~new_n9172_;
  assign new_n5699_ = ~new_n11405_;
  assign new_n11413_ = new_n9536_ & new_n9516_;
  assign new_n5700_ = ~new_n11413_;
  assign new_n11416_ = new_n7148_ & new_n11052_;
  assign new_n5701_ = ~new_n11416_;
  assign new_n11419_ = new_n11420_ & new_n11039_;
  assign new_n5702_ = ~new_n11419_;
  assign new_n11423_ = new_n9532_ & new_n9536_;
  assign new_n5703_ = ~new_n11423_;
  assign new_n11426_ = new_n11427_ & new_n9536_;
  assign new_n7370_ = ~new_n8774_;
  assign new_n5704_ = ~new_n11426_;
  assign new_n11430_ = new_n9536_ & new_n11431_;
  assign new_n5705_ = ~new_n11430_;
  assign new_n11470_ = IR_REG_26_ & new_n9536_;
  assign new_n5706_ = ~new_n11470_;
  assign new_n7577_ = new_n6002_ & new_n7579_;
  assign new_n5707_ = ~new_n7577_;
  assign new_n7583_ = new_n7584_ & new_n7585_;
  assign new_n5708_ = ~new_n7583_;
  assign new_n7598_ = new_n7599_ & new_n7600_;
  assign new_n7371_ = ~new_n9075_;
  assign new_n5709_ = ~new_n7598_;
  assign new_n7618_ = new_n6005_ & new_n7620_;
  assign new_n5710_ = ~new_n7618_;
  assign new_n7623_ = new_n7624_ & new_n7625_;
  assign new_n5711_ = ~new_n7623_;
  assign new_n7636_ = new_n7637_ & new_n5713_;
  assign new_n5712_ = ~new_n7636_;
  assign new_n7638_ = new_n7580_ & new_n7639_;
  assign new_n5713_ = ~new_n7638_;
  assign new_n7658_ = new_n6008_ & new_n5715_;
  assign new_n7372_ = ~new_n9060_;
  assign new_n5714_ = ~new_n7658_;
  assign new_n7660_ = new_n7586_ & new_n7661_;
  assign new_n5715_ = ~new_n7660_;
  assign new_n7665_ = new_n7666_ & new_n5717_;
  assign new_n5716_ = ~new_n7665_;
  assign new_n7667_ = new_n7668_ & new_n7580_;
  assign new_n5717_ = ~new_n7667_;
  assign new_n7679_ = new_n7680_ & new_n5719_;
  assign new_n5718_ = ~new_n7679_;
  assign new_n7681_ = new_n7682_ & new_n7580_;
  assign new_n7373_ = ~new_n9838_;
  assign new_n5719_ = ~new_n7681_;
  assign new_n7702_ = new_n6011_ & new_n5721_;
  assign new_n5720_ = ~new_n7702_;
  assign new_n7704_ = new_n7586_ & new_n7705_;
  assign new_n5721_ = ~new_n7704_;
  assign new_n7709_ = new_n7710_ & new_n5723_;
  assign new_n5722_ = ~new_n7709_;
  assign new_n7711_ = new_n7712_ & new_n7580_;
  assign new_n5723_ = ~new_n7711_;
  assign new_n7801_ = new_n6236_ | new_n6641_;
  assign new_n7374_ = ~new_n9612_;
  assign new_n5724_ = ~new_n7801_;
  assign new_n7821_ = new_n6238_ | new_n6643_;
  assign new_n5725_ = ~new_n7821_;
  assign new_n7838_ = new_n6240_ | new_n6645_;
  assign new_n5726_ = ~new_n7838_;
  assign new_n7855_ = new_n6242_ | new_n6647_;
  assign new_n5727_ = ~new_n7855_;
  assign new_n7872_ = new_n6244_ | new_n6649_;
  assign new_n5728_ = ~new_n7872_;
  assign new_n7889_ = new_n6246_ | new_n6651_;
  assign new_n7375_ = ~new_n9972_;
  assign new_n5729_ = ~new_n7889_;
  assign new_n7906_ = new_n6248_ | new_n6653_;
  assign new_n5730_ = ~new_n7906_;
  assign new_n7923_ = new_n6250_ | new_n6655_;
  assign new_n5731_ = ~new_n7923_;
  assign new_n7940_ = new_n6252_ | new_n6657_;
  assign new_n5732_ = ~new_n7940_;
  assign new_n7957_ = new_n6254_ | new_n6659_;
  assign new_n5733_ = ~new_n7957_;
  assign new_n7974_ = new_n6256_ | new_n6661_;
  assign new_n7376_ = ~new_n9597_;
  assign new_n5734_ = ~new_n7974_;
  assign new_n7991_ = new_n6258_ | new_n6663_;
  assign new_n5735_ = ~new_n7991_;
  assign new_n8008_ = new_n6260_ | new_n6665_;
  assign new_n5736_ = ~new_n8008_;
  assign new_n8025_ = new_n6262_ | new_n6667_;
  assign new_n5737_ = ~new_n8025_;
  assign new_n8042_ = new_n6264_ | new_n6669_;
  assign new_n5738_ = ~new_n8042_;
  assign new_n8059_ = new_n6266_ | new_n6671_;
  assign new_n7377_ = ~new_n10200_;
  assign new_n5739_ = ~new_n8059_;
  assign new_n8076_ = new_n6268_ | new_n6673_;
  assign new_n5740_ = ~new_n8076_;
  assign new_n8093_ = new_n6270_ | new_n6675_;
  assign new_n5741_ = ~new_n8093_;
  assign new_n8110_ = new_n6272_ | new_n6677_;
  assign new_n5742_ = ~new_n8110_;
  assign new_n8129_ = new_n6274_ | new_n6679_;
  assign new_n5743_ = ~new_n8129_;
  assign new_n8146_ = new_n6276_ | new_n6681_;
  assign new_n11172_ = new_n11398_ & REG1_REG_5_;
  assign new_n7378_ = ~new_n10070_;
  assign new_n5744_ = ~new_n8146_;
  assign new_n8164_ = new_n6278_ | new_n6683_;
  assign new_n5745_ = ~new_n8164_;
  assign new_n8181_ = new_n6280_ | new_n6685_;
  assign new_n5746_ = ~new_n8181_;
  assign new_n8199_ = new_n6282_ | new_n6687_;
  assign new_n5747_ = ~new_n8199_;
  assign new_n8216_ = new_n8217_ | new_n6689_;
  assign new_n5748_ = ~new_n8216_;
  assign new_n8232_ = new_n6285_ | new_n6691_;
  assign new_n7379_ = ~new_n8189_;
  assign new_n5749_ = ~new_n8232_;
  assign new_n8249_ = new_n6287_ | new_n6693_;
  assign new_n5750_ = ~new_n8249_;
  assign new_n8267_ = new_n6289_ | new_n6695_;
  assign new_n5751_ = ~new_n8267_;
  assign new_n8302_ = new_n8304_ & new_n7105_;
  assign new_n5752_ = ~new_n8302_;
  assign new_n8306_ = REG1_REG_30_ & new_n7564_;
  assign new_n5753_ = ~new_n8306_;
  assign new_n8309_ = REG1_REG_29_ & new_n7564_;
  assign new_n7380_ = ~new_n8119_;
  assign new_n5754_ = ~new_n8309_;
  assign new_n8312_ = REG1_REG_28_ & new_n7564_;
  assign new_n5755_ = ~new_n8312_;
  assign new_n8315_ = REG1_REG_27_ & new_n7564_;
  assign new_n5756_ = ~new_n8315_;
  assign new_n8318_ = REG1_REG_26_ & new_n7564_;
  assign new_n5757_ = ~new_n8318_;
  assign new_n8321_ = REG1_REG_25_ & new_n7564_;
  assign new_n5758_ = ~new_n8321_;
  assign new_n8324_ = REG1_REG_24_ & new_n7564_;
  assign new_n7381_ = ~new_n8015_;
  assign new_n5759_ = ~new_n8324_;
  assign new_n8327_ = REG1_REG_23_ & new_n7564_;
  assign new_n5760_ = ~new_n8327_;
  assign new_n8330_ = REG1_REG_22_ & new_n7564_;
  assign new_n5761_ = ~new_n8330_;
  assign new_n8333_ = REG1_REG_21_ & new_n7564_;
  assign new_n5762_ = ~new_n8333_;
  assign new_n8336_ = REG1_REG_20_ & new_n7564_;
  assign new_n5763_ = ~new_n8336_;
  assign new_n8339_ = REG1_REG_19_ & new_n7564_;
  assign new_n7382_ = ~new_n8049_;
  assign new_n5764_ = ~new_n8339_;
  assign new_n8342_ = REG1_REG_18_ & new_n7564_;
  assign new_n5765_ = ~new_n8342_;
  assign new_n8345_ = REG1_REG_17_ & new_n7564_;
  assign new_n5766_ = ~new_n8345_;
  assign new_n8348_ = REG1_REG_16_ & new_n7564_;
  assign new_n5767_ = ~new_n8348_;
  assign new_n8351_ = REG1_REG_15_ & new_n7564_;
  assign new_n5768_ = ~new_n8351_;
  assign new_n8354_ = REG1_REG_14_ & new_n7564_;
  assign new_n7383_ = ~new_n9927_;
  assign new_n5769_ = ~new_n8354_;
  assign new_n8357_ = REG1_REG_13_ & new_n7564_;
  assign new_n5770_ = ~new_n8357_;
  assign new_n8360_ = REG1_REG_12_ & new_n7564_;
  assign new_n5771_ = ~new_n8360_;
  assign new_n8363_ = REG1_REG_11_ & new_n7564_;
  assign new_n5772_ = ~new_n8363_;
  assign new_n8366_ = REG1_REG_10_ & new_n7564_;
  assign new_n5773_ = ~new_n8366_;
  assign new_n8369_ = REG1_REG_9_ & new_n7564_;
  assign new_n7384_ = ~new_n9868_;
  assign new_n5774_ = ~new_n8369_;
  assign new_n8372_ = REG1_REG_8_ & new_n7564_;
  assign new_n5775_ = ~new_n8372_;
  assign new_n8375_ = REG1_REG_7_ & new_n7564_;
  assign new_n5776_ = ~new_n8375_;
  assign new_n8378_ = REG1_REG_6_ & new_n7564_;
  assign new_n5777_ = ~new_n8378_;
  assign new_n8381_ = REG1_REG_5_ & new_n7564_;
  assign new_n5778_ = ~new_n8381_;
  assign new_n8384_ = REG1_REG_4_ & new_n7564_;
  assign new_n7947_ = DATAI_20_ & new_n7551_;
  assign new_n5779_ = ~new_n8384_;
  assign new_n8387_ = REG1_REG_3_ & new_n7564_;
  assign new_n5780_ = ~new_n8387_;
  assign new_n8390_ = REG1_REG_2_ & new_n7564_;
  assign new_n5781_ = ~new_n8390_;
  assign new_n8393_ = REG1_REG_1_ & new_n7564_;
  assign new_n5782_ = ~new_n8393_;
  assign new_n8396_ = REG1_REG_0_ & new_n7564_;
  assign new_n5783_ = ~new_n8396_;
  assign new_n8401_ = new_n8407_ & new_n7105_;
  assign new_n7385_ = ~new_n7947_;
  assign new_n5784_ = ~new_n8401_;
  assign new_n8409_ = new_n8407_ & new_n7106_;
  assign new_n5785_ = ~new_n8409_;
  assign new_n8421_ = new_n8407_ & new_n8310_;
  assign new_n5786_ = ~new_n8421_;
  assign new_n8458_ = new_n8407_ & new_n8313_;
  assign new_n5787_ = ~new_n8458_;
  assign new_n8484_ = new_n7828_ & new_n7361_;
  assign new_n5788_ = ~new_n8484_;
  assign new_n8487_ = new_n8407_ & new_n8316_;
  assign new_n7386_ = ~new_n8399_;
  assign new_n5789_ = ~new_n8487_;
  assign new_n8523_ = new_n8407_ & new_n8319_;
  assign new_n5790_ = ~new_n8523_;
  assign new_n8555_ = new_n8407_ & new_n8322_;
  assign new_n5791_ = ~new_n8555_;
  assign new_n8574_ = new_n8407_ & new_n8325_;
  assign new_n5792_ = ~new_n8574_;
  assign new_n8600_ = new_n8407_ & new_n8328_;
  assign new_n5793_ = ~new_n8600_;
  assign new_n8638_ = new_n7913_ & new_n7362_;
  assign new_n7061_ = ~new_n11172_;
  assign new_n7387_ = ~new_n10410_;
  assign new_n5794_ = ~new_n8638_;
  assign new_n8641_ = new_n8407_ & new_n8331_;
  assign new_n5795_ = ~new_n8641_;
  assign new_n8676_ = new_n8407_ & new_n8334_;
  assign new_n5796_ = ~new_n8676_;
  assign new_n8700_ = new_n8407_ & new_n8337_;
  assign new_n5797_ = ~new_n8700_;
  assign new_n8733_ = new_n8407_ & new_n8340_;
  assign new_n5798_ = ~new_n8733_;
  assign new_n8749_ = new_n7981_ & new_n8750_;
  assign new_n10410_ = new_n7393_ & new_n9043_;
  assign new_n5799_ = ~new_n8749_;
  assign new_n8752_ = new_n8407_ & new_n8343_;
  assign new_n5800_ = ~new_n8752_;
  assign new_n8773_ = new_n7370_ & new_n8775_;
  assign new_n5801_ = ~new_n8773_;
  assign new_n8779_ = new_n8407_ & new_n8346_;
  assign new_n5802_ = ~new_n8779_;
  assign new_n8807_ = new_n8407_ & new_n8349_;
  assign new_n5803_ = ~new_n8807_;
  assign new_n8844_ = new_n8407_ & new_n8352_;
  assign new_n7388_ = ~new_n10338_;
  assign new_n5804_ = ~new_n8844_;
  assign new_n8868_ = new_n8049_ & new_n8869_;
  assign new_n5805_ = ~new_n8868_;
  assign new_n8871_ = new_n8407_ & new_n8355_;
  assign new_n5806_ = ~new_n8871_;
  assign new_n8901_ = new_n8407_ & new_n8358_;
  assign new_n5807_ = ~new_n8901_;
  assign new_n8930_ = new_n8407_ & new_n8361_;
  assign new_n5808_ = ~new_n8930_;
  assign new_n8951_ = new_n8100_ & new_n8952_;
  assign new_n10338_ = new_n7480_ & new_n7407_;
  assign new_n5809_ = ~new_n8951_;
  assign new_n8954_ = new_n8407_ & new_n8364_;
  assign new_n5810_ = ~new_n8954_;
  assign new_n8983_ = new_n8984_ & new_n7124_;
  assign new_n5811_ = ~new_n8983_;
  assign new_n8991_ = new_n8407_ & new_n8367_;
  assign new_n5812_ = ~new_n8991_;
  assign new_n9027_ = new_n8407_ & new_n8370_;
  assign new_n5813_ = ~new_n9027_;
  assign new_n9042_ = new_n8154_ & new_n9043_;
  assign new_n7389_ = ~new_n10442_;
  assign new_n5814_ = ~new_n9042_;
  assign new_n9045_ = new_n8407_ & new_n8373_;
  assign new_n5815_ = ~new_n9045_;
  assign new_n9062_ = new_n9063_ & new_n7471_;
  assign new_n5816_ = ~new_n9062_;
  assign new_n9074_ = new_n7371_ & new_n9076_;
  assign new_n5817_ = ~new_n9074_;
  assign new_n9080_ = new_n8407_ & new_n8376_;
  assign new_n5818_ = ~new_n9080_;
  assign new_n9108_ = new_n8407_ & new_n8379_;
  assign new_n7390_ = ~new_n11106_;
  assign new_n5819_ = ~new_n9108_;
  assign new_n9123_ = new_n6113_ & new_n7520_;
  assign new_n5820_ = ~new_n9123_;
  assign new_n9143_ = new_n8407_ & new_n8382_;
  assign new_n5821_ = ~new_n9143_;
  assign new_n9175_ = new_n8407_ & new_n8385_;
  assign new_n5822_ = ~new_n9175_;
  assign new_n9198_ = new_n8407_ & new_n8388_;
  assign new_n5823_ = ~new_n9198_;
  assign new_n9215_ = new_n7257_ & new_n7442_;
  assign new_n7391_ = ~new_n8521_;
  assign new_n5824_ = ~new_n9215_;
  assign new_n9218_ = new_n8407_ & new_n8391_;
  assign new_n5825_ = ~new_n9218_;
  assign new_n9246_ = new_n8407_ & new_n8394_;
  assign new_n5826_ = ~new_n9246_;
  assign new_n9262_ = new_n8407_ & new_n7107_;
  assign new_n5827_ = ~new_n9262_;
  assign new_n9289_ = new_n7443_ & new_n5829_;
  assign new_n5828_ = ~new_n9289_;
  assign new_n9291_ = new_n7550_ & new_n7547_;
  assign new_n7392_ = ~new_n10445_;
  assign new_n5829_ = ~new_n9291_;
  assign new_n9295_ = new_n9293_ & new_n7108_;
  assign new_n5830_ = ~new_n9295_;
  assign new_n9298_ = D_REG_0_ & new_n7567_;
  assign new_n5831_ = ~new_n9298_;
  assign new_n9307_ = DATAI_30_ & n1332;
  assign new_n5832_ = ~new_n9307_;
  assign new_n9316_ = DATAI_29_ & n1332;
  assign new_n5833_ = ~new_n9316_;
  assign new_n9323_ = DATAI_28_ & n1332;
  assign new_n10445_ = new_n7815_ & new_n7461_;
  assign new_n5834_ = ~new_n9323_;
  assign new_n9327_ = new_n9313_ & new_n11447_;
  assign new_n5835_ = ~new_n9327_;
  assign new_n9331_ = DATAI_27_ & n1332;
  assign new_n5836_ = ~new_n9331_;
  assign new_n9335_ = new_n9313_ & new_n7481_;
  assign new_n5837_ = ~new_n9335_;
  assign new_n9340_ = DATAI_26_ & n1332;
  assign new_n5838_ = ~new_n9340_;
  assign new_n9345_ = DATAI_25_ & n1332;
  assign new_n7393_ = ~new_n8154_;
  assign new_n5839_ = ~new_n9345_;
  assign new_n9349_ = new_n9313_ & new_n9352_;
  assign new_n5840_ = ~new_n9349_;
  assign new_n9354_ = DATAI_24_ & n1332;
  assign new_n5841_ = ~new_n9354_;
  assign new_n9358_ = new_n9313_ & new_n7465_;
  assign new_n5842_ = ~new_n9358_;
  assign new_n9363_ = DATAI_23_ & n1332;
  assign new_n5843_ = ~new_n9363_;
  assign new_n9369_ = DATAI_22_ & n1332;
  assign new_n7062_ = ~new_n7591_;
  assign new_n7394_ = ~new_n9235_;
  assign new_n5844_ = ~new_n9369_;
  assign new_n9373_ = new_n9313_ & new_n7466_;
  assign new_n5845_ = ~new_n9373_;
  assign new_n9378_ = DATAI_21_ & n1332;
  assign new_n5846_ = ~new_n9378_;
  assign new_n9384_ = DATAI_20_ & n1332;
  assign new_n5847_ = ~new_n9384_;
  assign new_n9388_ = new_n9313_ & new_n7527_;
  assign new_n5848_ = ~new_n9388_;
  assign new_n9393_ = DATAI_19_ & n1332;
  assign new_n7913_ = DATAI_22_ & new_n7551_;
  assign new_n5849_ = ~new_n9393_;
  assign new_n9398_ = DATAI_18_ & n1332;
  assign new_n5850_ = ~new_n9398_;
  assign new_n9402_ = new_n9313_ & new_n7528_;
  assign new_n5851_ = ~new_n9402_;
  assign new_n9407_ = DATAI_17_ & n1332;
  assign new_n5852_ = ~new_n9407_;
  assign new_n9412_ = DATAI_16_ & n1332;
  assign new_n5853_ = ~new_n9412_;
  assign new_n9416_ = new_n9313_ & new_n7396_;
  assign new_n7395_ = ~new_n7913_;
  assign new_n5854_ = ~new_n9416_;
  assign new_n9421_ = DATAI_15_ & n1332;
  assign new_n5855_ = ~new_n9421_;
  assign new_n9427_ = DATAI_14_ & n1332;
  assign new_n5856_ = ~new_n9427_;
  assign new_n9431_ = new_n9313_ & new_n7397_;
  assign new_n5857_ = ~new_n9431_;
  assign new_n9436_ = DATAI_13_ & n1332;
  assign new_n5858_ = ~new_n9436_;
  assign new_n9442_ = DATAI_12_ & n1332;
  assign new_n7396_ = ~new_n9417_;
  assign new_n5859_ = ~new_n9442_;
  assign new_n9446_ = new_n9313_ & new_n7398_;
  assign new_n5860_ = ~new_n9446_;
  assign new_n9451_ = DATAI_11_ & n1332;
  assign new_n5861_ = ~new_n9451_;
  assign new_n9457_ = DATAI_10_ & n1332;
  assign new_n5862_ = ~new_n9457_;
  assign new_n9461_ = new_n9313_ & new_n7467_;
  assign new_n5863_ = ~new_n9461_;
  assign new_n9466_ = DATAI_9_ & n1332;
  assign new_n7397_ = ~new_n9432_;
  assign new_n5864_ = ~new_n9466_;
  assign new_n9472_ = DATAI_8_ & n1332;
  assign new_n5865_ = ~new_n9472_;
  assign new_n9476_ = new_n9313_ & new_n9484_;
  assign new_n5866_ = ~new_n9476_;
  assign new_n9480_ = DATAI_7_ & n1332;
  assign new_n5867_ = ~new_n9480_;
  assign new_n9487_ = DATAI_6_ & n1332;
  assign new_n5868_ = ~new_n9487_;
  assign new_n9491_ = new_n9313_ & new_n7468_;
  assign new_n7398_ = ~new_n9447_;
  assign new_n5869_ = ~new_n9491_;
  assign new_n9496_ = DATAI_5_ & n1332;
  assign new_n5870_ = ~new_n9496_;
  assign new_n9501_ = DATAI_4_ & n1332;
  assign new_n5871_ = ~new_n9501_;
  assign new_n9505_ = new_n9313_ & new_n7483_;
  assign new_n5872_ = ~new_n9505_;
  assign new_n9510_ = DATAI_3_ & n1332;
  assign new_n5873_ = ~new_n9510_;
  assign new_n9514_ = new_n9313_ & new_n9522_;
  assign new_n7399_ = ~new_n8967_;
  assign new_n5874_ = ~new_n9514_;
  assign new_n9518_ = DATAI_2_ & n1332;
  assign new_n5875_ = ~new_n9518_;
  assign new_n9525_ = DATAI_1_ & n1332;
  assign new_n5876_ = ~new_n9525_;
  assign new_n9529_ = new_n9313_ & new_n9530_;
  assign new_n5877_ = ~new_n9529_;
  assign new_n9534_ = IR_REG_0_ & new_n5879_;
  assign new_n5878_ = ~new_n9534_;
  assign new_n9535_ = new_n7553_ & new_n7552_;
  assign new_n7400_ = ~new_n9944_;
  assign new_n5879_ = ~new_n9535_;
  assign new_n9559_ = new_n7305_ & new_n7280_;
  assign new_n5880_ = ~new_n9559_;
  assign new_n10046_ = new_n9661_ & new_n9660_;
  assign new_n5881_ = ~new_n10046_;
  assign new_n10153_ = new_n6146_ & new_n7405_;
  assign new_n5882_ = ~new_n10153_;
  assign new_n10161_ = new_n7291_ & new_n5884_;
  assign new_n5883_ = ~new_n10161_;
  assign new_n10162_ = new_n9948_ & new_n7271_;
  assign new_n7401_ = ~new_n9352_;
  assign new_n5884_ = ~new_n10162_;
  assign new_n10168_ = new_n9865_ & new_n7384_;
  assign new_n5885_ = ~new_n10168_;
  assign new_n10180_ = new_n9852_ & new_n9851_;
  assign new_n5886_ = ~new_n10180_;
  assign new_n10226_ = new_n7412_ & new_n7305_;
  assign new_n5887_ = ~new_n10226_;
  assign new_n10287_ = new_n6148_ & new_n5889_;
  assign new_n5888_ = ~new_n10287_;
  assign new_n10289_ = new_n10290_ | new_n10291_;
  assign new_n9352_ = new_n7465_ & new_n9361_;
  assign new_n5889_ = ~new_n10289_;
  assign new_n10293_ = new_n6149_ & new_n5891_;
  assign new_n5890_ = ~new_n10293_;
  assign new_n10295_ = new_n10296_ | new_n10297_;
  assign new_n5891_ = ~new_n10295_;
  assign new_n10302_ = new_n6150_ & new_n5893_;
  assign new_n5892_ = ~new_n10302_;
  assign new_n10304_ = new_n10305_ | new_n10306_;
  assign new_n5893_ = ~new_n10304_;
  assign new_n10309_ = new_n6151_ & new_n5895_;
  assign new_n9823_ = new_n10053_ & new_n10054_;
  assign new_n7402_ = ~new_n11179_;
  assign new_n5894_ = ~new_n10309_;
  assign new_n10311_ = new_n10312_ | new_n10313_;
  assign new_n5895_ = ~new_n10311_;
  assign new_n10326_ = new_n10704_ & new_n5897_;
  assign new_n5896_ = ~new_n10326_;
  assign new_n10327_ = new_n6156_ & new_n10329_;
  assign new_n5897_ = ~new_n10327_;
  assign new_n10341_ = new_n10342_ & new_n5899_;
  assign new_n5898_ = ~new_n10341_;
  assign new_n10343_ = new_n10344_ & new_n5900_;
  assign new_n7403_ = ~new_n9059_;
  assign new_n5899_ = ~new_n10343_;
  assign new_n10345_ = new_n10346_ & new_n5901_;
  assign new_n5900_ = ~new_n10345_;
  assign new_n10347_ = new_n10348_ & new_n5902_;
  assign new_n5901_ = ~new_n10347_;
  assign new_n10349_ = new_n10350_ & new_n5903_;
  assign new_n5902_ = ~new_n10349_;
  assign new_n10351_ = new_n10352_ & new_n5904_;
  assign new_n5903_ = ~new_n10351_;
  assign new_n10353_ = new_n8621_ & new_n5905_;
  assign new_n9522_ = new_n11428_ & new_n11427_;
  assign new_n5904_ = ~new_n10353_;
  assign new_n10354_ = new_n10355_ & new_n5906_;
  assign new_n5905_ = ~new_n10354_;
  assign new_n10356_ = new_n10357_ & new_n5907_;
  assign new_n5906_ = ~new_n10356_;
  assign new_n10358_ = new_n10359_ & new_n5908_;
  assign new_n5907_ = ~new_n10358_;
  assign new_n10360_ = new_n10361_ & new_n5909_;
  assign new_n5908_ = ~new_n10360_;
  assign new_n10362_ = new_n10363_ & new_n5910_;
  assign new_n7404_ = ~new_n9522_;
  assign new_n5909_ = ~new_n10362_;
  assign new_n10364_ = new_n10365_ & new_n5911_;
  assign new_n5910_ = ~new_n10364_;
  assign new_n10366_ = new_n10367_ & new_n5912_;
  assign new_n5911_ = ~new_n10366_;
  assign new_n10368_ = new_n10369_ & new_n10370_;
  assign new_n5912_ = ~new_n10368_;
  assign new_n10394_ = new_n6154_ & new_n7473_;
  assign new_n5913_ = ~new_n10394_;
  assign new_n10475_ = new_n7524_ & new_n5915_;
  assign new_n9761_ = new_n10155_ & new_n10156_;
  assign new_n5914_ = ~new_n10475_;
  assign new_n10476_ = new_n8468_ & new_n7539_;
  assign new_n5915_ = ~new_n10476_;
  assign new_n10485_ = new_n8472_ | new_n6711_;
  assign new_n5916_ = ~new_n10485_;
  assign new_n10532_ = new_n7418_ & new_n5918_;
  assign new_n5917_ = ~new_n10532_;
  assign new_n10533_ = new_n9280_ & new_n7701_;
  assign new_n5918_ = ~new_n10533_;
  assign new_n10545_ = new_n7135_ & new_n5920_;
  assign new_n7405_ = ~new_n9761_;
  assign new_n5919_ = ~new_n10545_;
  assign new_n10547_ = new_n7459_ & new_n5921_;
  assign new_n5920_ = ~new_n10547_;
  assign new_n10548_ = new_n6162_ & new_n7525_;
  assign new_n5921_ = ~new_n10548_;
  assign new_n10557_ = new_n9059_ & new_n7387_;
  assign new_n5922_ = ~new_n10557_;
  assign new_n10560_ = new_n9122_ & new_n7473_;
  assign new_n5923_ = ~new_n10560_;
  assign new_n10571_ = new_n6164_ & new_n7542_;
  assign new_n7406_ = ~new_n10415_;
  assign new_n5924_ = ~new_n10571_;
  assign new_n10576_ = new_n7409_ & new_n5926_;
  assign new_n5925_ = ~new_n10576_;
  assign new_n10577_ = new_n10411_ & new_n7523_;
  assign new_n5926_ = ~new_n10577_;
  assign new_n10581_ = new_n6304_ | new_n6714_;
  assign new_n5927_ = ~new_n10581_;
  assign new_n10624_ = new_n7543_ & new_n10625_;
  assign new_n5928_ = ~new_n10624_;
  assign new_n10645_ = new_n7458_ & new_n5930_;
  assign new_n8416_ = DATAI_30_ & new_n7551_;
  assign new_n5929_ = ~new_n10645_;
  assign new_n10646_ = new_n8968_ & new_n7281_;
  assign new_n5930_ = ~new_n10646_;
  assign new_n5931_ = ~new_n9424_;
  assign new_n5932_ = ~new_n9439_;
  assign new_n10706_ = n1341 & new_n7521_;
  assign new_n5933_ = ~new_n10706_;
  assign new_n10716_ = n1341 & new_n7480_;
  assign new_n5934_ = ~new_n10716_;
  assign new_n10722_ = n1341 & new_n7815_;
  assign new_n7407_ = ~new_n8416_;
  assign new_n5935_ = ~new_n10722_;
  assign new_n10732_ = n1341 & new_n8454_;
  assign new_n5936_ = ~new_n10732_;
  assign new_n10742_ = n1341 & new_n8483_;
  assign new_n5937_ = ~new_n10742_;
  assign new_n10750_ = n1341 & new_n8553_;
  assign new_n5938_ = ~new_n10750_;
  assign new_n10763_ = n1341 & new_n8552_;
  assign new_n5939_ = ~new_n10763_;
  assign new_n10771_ = n1341 & new_n8521_;
  assign new_n7408_ = ~new_n10416_;
  assign new_n5940_ = ~new_n10771_;
  assign new_n10784_ = n1341 & new_n8596_;
  assign new_n5941_ = ~new_n10784_;
  assign new_n10792_ = n1341 & new_n8637_;
  assign new_n5942_ = ~new_n10792_;
  assign new_n10803_ = n1341 & new_n8674_;
  assign new_n5943_ = ~new_n10803_;
  assign new_n10812_ = n1341 & new_n8728_;
  assign new_n5944_ = ~new_n10812_;
  assign new_n10824_ = n1341 & new_n8729_;
  assign new_n7063_ = ~new_n9823_;
  assign new_n7409_ = ~new_n10414_;
  assign new_n5945_ = ~new_n10824_;
  assign new_n10832_ = n1341 & new_n8750_;
  assign new_n5946_ = ~new_n10832_;
  assign new_n10845_ = n1341 & new_n8774_;
  assign new_n5947_ = ~new_n10845_;
  assign new_n10853_ = n1341 & new_n8805_;
  assign new_n5948_ = ~new_n10853_;
  assign new_n10866_ = n1341 & new_n8841_;
  assign new_n5949_ = ~new_n10866_;
  assign new_n10874_ = n1341 & new_n8869_;
  assign new_n7410_ = ~new_n9300_;
  assign new_n5950_ = ~new_n10874_;
  assign new_n10886_ = n1341 & new_n8927_;
  assign new_n5951_ = ~new_n10886_;
  assign new_n10894_ = n1341 & new_n8928_;
  assign new_n5952_ = ~new_n10894_;
  assign new_n10907_ = n1341 & new_n8952_;
  assign new_n5953_ = ~new_n10907_;
  assign new_n10915_ = n1341 & new_n9024_;
  assign new_n5954_ = ~new_n10915_;
  assign new_n10928_ = n1341 & new_n9025_;
  assign new_n7411_ = ~new_n8290_;
  assign new_n5955_ = ~new_n10928_;
  assign new_n10936_ = n1341 & new_n9043_;
  assign new_n5956_ = ~new_n10936_;
  assign new_n10949_ = n1341 & new_n9075_;
  assign new_n5957_ = ~new_n10949_;
  assign new_n10958_ = n1341 & new_n9106_;
  assign new_n5958_ = ~new_n10958_;
  assign new_n10968_ = n1341 & new_n9173_;
  assign new_n5959_ = ~new_n10968_;
  assign new_n10976_ = n1341 & new_n9171_;
  assign new_n7412_ = ~new_n9563_;
  assign new_n5960_ = ~new_n10976_;
  assign new_n10985_ = n1341 & new_n8262_;
  assign new_n5961_ = ~new_n10985_;
  assign new_n10993_ = n1341 & new_n9216_;
  assign new_n5962_ = ~new_n10993_;
  assign new_n11001_ = n1341 & new_n10442_;
  assign new_n5963_ = ~new_n11001_;
  assign new_n11009_ = n1341 & new_n10586_;
  assign new_n5964_ = ~new_n11009_;
  assign new_n11046_ = new_n6203_ & new_n5966_;
  assign new_n10419_ = new_n8483_ & new_n7457_;
  assign new_n5965_ = ~new_n11046_;
  assign new_n11048_ = new_n7586_ & new_n11049_;
  assign new_n5966_ = ~new_n11048_;
  assign new_n11053_ = new_n11054_ & new_n5968_;
  assign new_n5967_ = ~new_n11053_;
  assign new_n11055_ = new_n11056_ & new_n7580_;
  assign new_n5968_ = ~new_n11055_;
  assign new_n11067_ = new_n11068_ & new_n5970_;
  assign new_n5969_ = ~new_n11067_;
  assign new_n11069_ = new_n7580_ & new_n7192_;
  assign new_n7413_ = ~new_n10419_;
  assign new_n5970_ = ~new_n11069_;
  assign new_n11086_ = new_n11087_ & new_n5972_;
  assign new_n5971_ = ~new_n11086_;
  assign new_n11088_ = new_n7580_ & new_n11089_;
  assign new_n5972_ = ~new_n11088_;
  assign new_n11160_ = new_n11161_ & new_n5974_;
  assign new_n5973_ = ~new_n11160_;
  assign new_n11162_ = new_n7580_ & new_n7193_;
  assign new_n5974_ = ~new_n11162_;
  assign new_n11168_ = new_n6211_ & new_n11170_;
  assign new_n7414_ = ~new_n10409_;
  assign new_n5975_ = ~new_n11168_;
  assign new_n11180_ = new_n11181_ & new_n5977_;
  assign new_n5976_ = ~new_n11180_;
  assign new_n11182_ = new_n7580_ & new_n11183_;
  assign new_n5977_ = ~new_n11182_;
  assign new_n11200_ = new_n6214_ & new_n5979_;
  assign new_n5978_ = ~new_n11200_;
  assign new_n11202_ = new_n7586_ & new_n11203_;
  assign new_n5979_ = ~new_n11202_;
  assign new_n11207_ = new_n11208_ & new_n5981_;
  assign new_n10409_ = new_n7442_ & new_n9216_;
  assign new_n5980_ = ~new_n11207_;
  assign new_n11209_ = new_n11210_ & new_n7580_;
  assign new_n5981_ = ~new_n11209_;
  assign new_n11219_ = new_n11220_ & new_n5983_;
  assign new_n5982_ = ~new_n11219_;
  assign new_n11221_ = new_n7580_ & new_n7194_;
  assign new_n5983_ = ~new_n11221_;
  assign new_n11238_ = new_n6217_ & new_n5985_;
  assign new_n5984_ = ~new_n11238_;
  assign new_n11240_ = new_n7586_ & new_n11241_;
  assign new_n7415_ = ~new_n9005_;
  assign new_n5985_ = ~new_n11240_;
  assign new_n11244_ = new_n11245_ & new_n5987_;
  assign new_n5986_ = ~new_n11244_;
  assign new_n11246_ = new_n7580_ & new_n11247_;
  assign new_n5987_ = ~new_n11246_;
  assign new_n11257_ = new_n11258_ & new_n5989_;
  assign new_n5988_ = ~new_n11257_;
  assign new_n11259_ = new_n7580_ & new_n7195_;
  assign new_n5989_ = ~new_n11259_;
  assign new_n11276_ = new_n6220_ & new_n5991_;
  assign new_n7416_ = ~new_n9762_;
  assign new_n5990_ = ~new_n11276_;
  assign new_n11278_ = new_n7586_ & new_n11279_;
  assign new_n5991_ = ~new_n11278_;
  assign new_n11284_ = new_n11285_ & new_n5993_;
  assign new_n5992_ = ~new_n11284_;
  assign new_n11286_ = new_n7580_ & new_n11287_;
  assign new_n5993_ = ~new_n11286_;
  assign new_n11297_ = new_n11298_ & new_n5995_;
  assign new_n5994_ = ~new_n11297_;
  assign new_n11299_ = new_n11300_ & new_n7580_;
  assign new_n9693_ = new_n10094_ & new_n10095_;
  assign new_n7417_ = ~new_n10452_;
  assign new_n5995_ = ~new_n11299_;
  assign new_n5996_ = ~new_n9454_;
  assign new_n11367_ = new_n9462_ & new_n7163_;
  assign new_n5997_ = ~new_n11367_;
  assign new_n5998_ = ~new_n9521_;
  assign new_n5999_ = ~new_n9483_;
  assign new_n11440_ = new_n9374_ & new_n7164_;
  assign new_n6000_ = ~new_n11440_;
  assign new_n11458_ = new_n9359_ & new_n7165_;
  assign new_n6001_ = ~new_n11458_;
  assign new_n7418_ = ~new_n8300_;
  assign new_n7578_ = new_n7586_ & new_n7582_;
  assign new_n6002_ = ~new_n7578_;
  assign new_n7604_ = new_n6004_ & new_n7607_;
  assign new_n6003_ = ~new_n7604_;
  assign new_n7606_ = new_n7586_ & new_n7601_;
  assign new_n6004_ = ~new_n7606_;
  assign new_n7619_ = new_n7586_ & new_n7622_;
  assign new_n6005_ = ~new_n7619_;
  assign new_n6006_ = ~new_n7645_;
  assign new_n7647_ = new_n7650_ & new_n7580_;
  assign new_n8776_ = new_n8015_ & new_n8805_;
  assign new_n6007_ = ~new_n7647_;
  assign new_n7659_ = new_n7580_ & new_n7663_;
  assign new_n6008_ = ~new_n7659_;
  assign new_n6009_ = ~new_n7690_;
  assign new_n7691_ = new_n7580_ & new_n7694_;
  assign new_n6010_ = ~new_n7691_;
  assign new_n7703_ = new_n7580_ & new_n7707_;
  assign new_n6011_ = ~new_n7703_;
  assign new_n7721_ = new_n7646_ & new_n7003_;
  assign new_n6012_ = ~new_n7721_;
  assign new_n7419_ = ~new_n8776_;
  assign new_n7800_ = new_n6237_ | new_n6642_;
  assign new_n6013_ = ~new_n7800_;
  assign new_n7820_ = new_n6239_ | new_n6644_;
  assign new_n6014_ = ~new_n7820_;
  assign new_n7837_ = new_n6241_ | new_n6646_;
  assign new_n6015_ = ~new_n7837_;
  assign new_n7854_ = new_n6243_ | new_n6648_;
  assign new_n6016_ = ~new_n7854_;
  assign new_n7871_ = new_n6245_ | new_n6650_;
  assign new_n6017_ = ~new_n7871_;
  assign new_n9077_ = new_n8189_ & new_n9106_;
  assign new_n7888_ = new_n6247_ | new_n6652_;
  assign new_n6018_ = ~new_n7888_;
  assign new_n7905_ = new_n6249_ | new_n6654_;
  assign new_n6019_ = ~new_n7905_;
  assign new_n7922_ = new_n6251_ | new_n6656_;
  assign new_n6020_ = ~new_n7922_;
  assign new_n7939_ = new_n6253_ | new_n6658_;
  assign new_n6021_ = ~new_n7939_;
  assign new_n7956_ = new_n6255_ | new_n6660_;
  assign new_n6022_ = ~new_n7956_;
  assign new_n7420_ = ~new_n9077_;
  assign new_n7973_ = new_n6257_ | new_n6662_;
  assign new_n6023_ = ~new_n7973_;
  assign new_n7990_ = new_n6259_ | new_n6664_;
  assign new_n6024_ = ~new_n7990_;
  assign new_n8007_ = new_n6261_ | new_n6666_;
  assign new_n6025_ = ~new_n8007_;
  assign new_n8024_ = new_n6263_ | new_n6668_;
  assign new_n6026_ = ~new_n8024_;
  assign new_n8041_ = new_n6265_ | new_n6670_;
  assign new_n6027_ = ~new_n8041_;
  assign new_n9141_ = new_n9172_ & new_n9171_;
  assign new_n8058_ = new_n6267_ | new_n6672_;
  assign new_n6028_ = ~new_n8058_;
  assign new_n8075_ = new_n6269_ | new_n6674_;
  assign new_n6029_ = ~new_n8075_;
  assign new_n8092_ = new_n6271_ | new_n6676_;
  assign new_n6030_ = ~new_n8092_;
  assign new_n8109_ = new_n6273_ | new_n6678_;
  assign new_n6031_ = ~new_n8109_;
  assign new_n8128_ = new_n6275_ | new_n6680_;
  assign new_n6032_ = ~new_n8128_;
  assign new_n7421_ = ~new_n9141_;
  assign new_n8145_ = new_n6277_ | new_n6682_;
  assign new_n6033_ = ~new_n8145_;
  assign new_n8163_ = new_n6279_ | new_n6684_;
  assign new_n6034_ = ~new_n8163_;
  assign new_n8180_ = new_n6281_ | new_n6686_;
  assign new_n6035_ = ~new_n8180_;
  assign new_n8198_ = new_n6283_ | new_n6688_;
  assign new_n6036_ = ~new_n8198_;
  assign new_n8215_ = new_n6284_ | new_n6690_;
  assign new_n6037_ = ~new_n8215_;
  assign new_n10418_ = new_n8521_ & new_n7454_;
  assign new_n8231_ = new_n6286_ | new_n6692_;
  assign new_n6038_ = ~new_n8231_;
  assign new_n8248_ = new_n6288_ | new_n6694_;
  assign new_n6039_ = ~new_n8248_;
  assign new_n8266_ = new_n6290_ | new_n6696_;
  assign new_n6040_ = ~new_n8266_;
  assign new_n8301_ = REG1_REG_31_ & new_n7564_;
  assign new_n6041_ = ~new_n8301_;
  assign new_n8305_ = new_n8304_ & new_n7106_;
  assign new_n6042_ = ~new_n8305_;
  assign new_n7422_ = ~new_n10418_;
  assign new_n8308_ = new_n8304_ & new_n8310_;
  assign new_n6043_ = ~new_n8308_;
  assign new_n8311_ = new_n8304_ & new_n8313_;
  assign new_n6044_ = ~new_n8311_;
  assign new_n8314_ = new_n8304_ & new_n8316_;
  assign new_n6045_ = ~new_n8314_;
  assign new_n8317_ = new_n8304_ & new_n8319_;
  assign new_n6046_ = ~new_n8317_;
  assign new_n8320_ = new_n8304_ & new_n8322_;
  assign new_n6047_ = ~new_n8320_;
  assign new_n7064_ = ~new_n9693_;
  assign new_n7423_ = ~new_n9554_;
  assign new_n8323_ = new_n8304_ & new_n8325_;
  assign new_n6048_ = ~new_n8323_;
  assign new_n8326_ = new_n8304_ & new_n8328_;
  assign new_n6049_ = ~new_n8326_;
  assign new_n8329_ = new_n8304_ & new_n8331_;
  assign new_n6050_ = ~new_n8329_;
  assign new_n8332_ = new_n8304_ & new_n8334_;
  assign new_n6051_ = ~new_n8332_;
  assign new_n8335_ = new_n8304_ & new_n8337_;
  assign new_n6052_ = ~new_n8335_;
  assign new_n7424_ = ~new_n11136_;
  assign new_n8338_ = new_n8304_ & new_n8340_;
  assign new_n6053_ = ~new_n8338_;
  assign new_n8341_ = new_n8304_ & new_n8343_;
  assign new_n6054_ = ~new_n8341_;
  assign new_n8344_ = new_n8304_ & new_n8346_;
  assign new_n6055_ = ~new_n8344_;
  assign new_n8347_ = new_n8304_ & new_n8349_;
  assign new_n6056_ = ~new_n8347_;
  assign new_n8350_ = new_n8304_ & new_n8352_;
  assign new_n6057_ = ~new_n8350_;
  assign new_n9185_ = new_n7525_ & new_n7459_;
  assign new_n8353_ = new_n8304_ & new_n8355_;
  assign new_n6058_ = ~new_n8353_;
  assign new_n8356_ = new_n8304_ & new_n8358_;
  assign new_n6059_ = ~new_n8356_;
  assign new_n8359_ = new_n8304_ & new_n8361_;
  assign new_n6060_ = ~new_n8359_;
  assign new_n8362_ = new_n8304_ & new_n8364_;
  assign new_n6061_ = ~new_n8362_;
  assign new_n8365_ = new_n8304_ & new_n8367_;
  assign new_n6062_ = ~new_n8365_;
  assign new_n7425_ = ~new_n9185_;
  assign new_n8368_ = new_n8304_ & new_n8370_;
  assign new_n6063_ = ~new_n8368_;
  assign new_n8371_ = new_n8304_ & new_n8373_;
  assign new_n6064_ = ~new_n8371_;
  assign new_n8374_ = new_n8304_ & new_n8376_;
  assign new_n6065_ = ~new_n8374_;
  assign new_n8377_ = new_n8304_ & new_n8379_;
  assign new_n6066_ = ~new_n8377_;
  assign new_n8380_ = new_n8304_ & new_n8382_;
  assign new_n6067_ = ~new_n8380_;
  assign new_n7426_ = ~new_n11036_;
  assign new_n8383_ = new_n8304_ & new_n8385_;
  assign new_n6068_ = ~new_n8383_;
  assign new_n8386_ = new_n8304_ & new_n8388_;
  assign new_n6069_ = ~new_n8386_;
  assign new_n8389_ = new_n8304_ & new_n8391_;
  assign new_n6070_ = ~new_n8389_;
  assign new_n8392_ = new_n8304_ & new_n8394_;
  assign new_n6071_ = ~new_n8392_;
  assign new_n8395_ = new_n8304_ & new_n7107_;
  assign new_n6072_ = ~new_n8395_;
  assign new_n7427_ = ~new_n9256_;
  assign new_n8400_ = REG0_REG_31_ & new_n7565_;
  assign new_n6073_ = ~new_n8400_;
  assign new_n8408_ = REG0_REG_30_ & new_n7565_;
  assign new_n6074_ = ~new_n8408_;
  assign new_n8436_ = new_n6291_ | new_n6699_;
  assign new_n6075_ = ~new_n8436_;
  assign new_n8420_ = REG0_REG_29_ & new_n7565_;
  assign new_n6076_ = ~new_n8420_;
  assign new_n8457_ = REG0_REG_28_ & new_n7565_;
  assign new_n6077_ = ~new_n8457_;
  assign new_n7428_ = ~new_n9036_;
  assign new_n8514_ = new_n8516_ & new_n7298_;
  assign new_n6078_ = ~new_n8514_;
  assign new_n8486_ = REG0_REG_27_ & new_n7565_;
  assign new_n6079_ = ~new_n8486_;
  assign new_n8522_ = REG0_REG_26_ & new_n7565_;
  assign new_n6080_ = ~new_n8522_;
  assign new_n8571_ = new_n7879_ & new_n8521_;
  assign new_n6081_ = ~new_n8571_;
  assign new_n8554_ = REG0_REG_25_ & new_n7565_;
  assign new_n6082_ = ~new_n8554_;
  assign new_n7429_ = ~new_n9133_;
  assign new_n8573_ = REG0_REG_24_ & new_n7565_;
  assign new_n6083_ = ~new_n8573_;
  assign new_n6084_ = ~new_n8613_;
  assign new_n8599_ = REG0_REG_23_ & new_n7565_;
  assign new_n6085_ = ~new_n8599_;
  assign new_n8640_ = REG0_REG_22_ & new_n7565_;
  assign new_n6086_ = ~new_n8640_;
  assign new_n6087_ = ~new_n8693_;
  assign new_n8675_ = REG0_REG_21_ & new_n7565_;
  assign new_n6088_ = ~new_n8675_;
  assign new_n7430_ = ~new_n10882_;
  assign new_n8699_ = REG0_REG_20_ & new_n7565_;
  assign new_n6089_ = ~new_n8699_;
  assign new_n8732_ = REG0_REG_19_ & new_n7565_;
  assign new_n6090_ = ~new_n8732_;
  assign new_n8772_ = new_n7536_ & new_n7419_;
  assign new_n6091_ = ~new_n8772_;
  assign new_n8751_ = REG0_REG_18_ & new_n7565_;
  assign new_n6092_ = ~new_n8751_;
  assign new_n8778_ = REG0_REG_17_ & new_n7565_;
  assign new_n6093_ = ~new_n8778_;
  assign new_n10882_ = new_n10902_ & REG3_REG_12_;
  assign new_n8819_ = new_n7541_ & new_n7020_;
  assign new_n6094_ = ~new_n8819_;
  assign new_n8823_ = new_n6096_ & new_n7541_;
  assign new_n6095_ = ~new_n8823_;
  assign new_n8825_ = new_n8822_ & new_n7542_;
  assign new_n6096_ = ~new_n8825_;
  assign new_n8842_ = new_n7532_ & new_n7311_;
  assign new_n6097_ = ~new_n8842_;
  assign new_n8806_ = REG0_REG_16_ & new_n7565_;
  assign new_n6098_ = ~new_n8806_;
  assign new_n9244_ = new_n7389_ & new_n7549_;
  assign new_n8404_ = DATAI_31_ & new_n7551_;
  assign new_n8843_ = REG0_REG_15_ & new_n7565_;
  assign new_n6099_ = ~new_n8843_;
  assign new_n8870_ = REG0_REG_14_ & new_n7565_;
  assign new_n6100_ = ~new_n8870_;
  assign new_n8900_ = REG0_REG_13_ & new_n7565_;
  assign new_n6101_ = ~new_n8900_;
  assign new_n8929_ = REG0_REG_12_ & new_n7565_;
  assign new_n6102_ = ~new_n8929_;
  assign new_n8966_ = new_n7453_ & new_n7253_;
  assign new_n6103_ = ~new_n8966_;
  assign new_n7431_ = ~new_n8404_;
  assign new_n8970_ = new_n7211_ & new_n7453_;
  assign new_n6104_ = ~new_n8970_;
  assign new_n8953_ = REG0_REG_11_ & new_n7565_;
  assign new_n6105_ = ~new_n8953_;
  assign new_n9000_ = new_n7275_ & new_n7253_;
  assign new_n6106_ = ~new_n9000_;
  assign new_n8990_ = REG0_REG_10_ & new_n7565_;
  assign new_n6107_ = ~new_n8990_;
  assign new_n9026_ = REG0_REG_9_ & new_n7565_;
  assign new_n6108_ = ~new_n9026_;
  assign new_n11022_ = REG1_REG_0_ & IR_REG_0_;
  assign new_n9058_ = new_n7372_ & new_n7471_;
  assign new_n6109_ = ~new_n9058_;
  assign new_n9073_ = new_n7534_ & new_n7420_;
  assign new_n6110_ = ~new_n9073_;
  assign new_n9044_ = REG0_REG_8_ & new_n7565_;
  assign new_n6111_ = ~new_n9044_;
  assign new_n9079_ = REG0_REG_7_ & new_n7565_;
  assign new_n6112_ = ~new_n9079_;
  assign new_n9124_ = new_n7508_ & new_n7254_;
  assign new_n6113_ = ~new_n9124_;
  assign new_n7432_ = ~new_n11022_;
  assign new_n9107_ = REG0_REG_6_ & new_n7565_;
  assign new_n6114_ = ~new_n9107_;
  assign new_n9152_ = new_n7053_ & new_n7254_;
  assign new_n6115_ = ~new_n9152_;
  assign new_n9142_ = REG0_REG_5_ & new_n7565_;
  assign new_n6116_ = ~new_n9142_;
  assign new_n9174_ = REG0_REG_4_ & new_n7565_;
  assign new_n6117_ = ~new_n9174_;
  assign new_n9197_ = REG0_REG_3_ & new_n7565_;
  assign new_n6118_ = ~new_n9197_;
  assign new_n7433_ = ~new_n9020_;
  assign new_n9217_ = REG0_REG_2_ & new_n7565_;
  assign new_n6119_ = ~new_n9217_;
  assign new_n9245_ = REG0_REG_1_ & new_n7565_;
  assign new_n6120_ = ~new_n9245_;
  assign new_n9270_ = new_n6122_ & new_n8291_;
  assign new_n6121_ = ~new_n9270_;
  assign new_n9271_ = new_n8292_ | new_n8450_;
  assign new_n6122_ = ~new_n9271_;
  assign new_n9261_ = REG0_REG_0_ & new_n7565_;
  assign new_n6123_ = ~new_n9261_;
  assign new_n7434_ = ~new_n8614_;
  assign new_n9288_ = new_n10324_ | new_n9292_;
  assign new_n6124_ = ~new_n9288_;
  assign new_n9294_ = D_REG_1_ & new_n7567_;
  assign new_n6125_ = ~new_n9294_;
  assign new_n9297_ = new_n9293_ & new_n7076_;
  assign new_n6126_ = ~new_n9297_;
  assign new_n9301_ = DATAI_31_ & n1332;
  assign new_n6127_ = ~new_n9301_;
  assign new_n9328_ = new_n7552_ | new_n11447_;
  assign new_n6128_ = ~new_n9328_;
  assign new_n7435_ = ~new_n8471_;
  assign new_n9337_ = new_n7481_ | new_n7552_;
  assign new_n6129_ = ~new_n9337_;
  assign new_n9360_ = new_n7552_ | new_n7465_;
  assign new_n6130_ = ~new_n9360_;
  assign new_n9375_ = new_n7552_ | new_n7466_;
  assign new_n6131_ = ~new_n9375_;
  assign new_n9390_ = new_n7527_ | new_n7552_;
  assign new_n6132_ = ~new_n9390_;
  assign new_n9404_ = new_n7528_ | new_n7552_;
  assign new_n6133_ = ~new_n9404_;
  assign new_n7436_ = ~new_n8923_;
  assign new_n9418_ = new_n7552_ | new_n7396_;
  assign new_n6134_ = ~new_n9418_;
  assign new_n9433_ = new_n7552_ | new_n7397_;
  assign new_n6135_ = ~new_n9433_;
  assign new_n9448_ = new_n7552_ | new_n7398_;
  assign new_n6136_ = ~new_n9448_;
  assign new_n9463_ = new_n7552_ | new_n7467_;
  assign new_n6137_ = ~new_n9463_;
  assign new_n9477_ = new_n7552_ | new_n9484_;
  assign new_n6138_ = ~new_n9477_;
  assign new_n7437_ = ~new_n8066_;
  assign new_n9493_ = new_n7552_ | new_n7468_;
  assign new_n6139_ = ~new_n9493_;
  assign new_n9507_ = new_n7552_ | new_n7483_;
  assign new_n6140_ = ~new_n9507_;
  assign new_n9515_ = new_n7552_ | new_n9522_;
  assign new_n6141_ = ~new_n9515_;
  assign new_n9531_ = new_n7552_ | new_n9530_;
  assign new_n6142_ = ~new_n9531_;
  assign new_n9533_ = DATAI_0_ & n1332;
  assign new_n6143_ = ~new_n9533_;
  assign new_n7438_ = ~new_n7964_;
  assign new_n10067_ = new_n10069_ & new_n7378_;
  assign new_n6144_ = ~new_n10067_;
  assign new_n10136_ = new_n10137_ & new_n7263_;
  assign new_n6145_ = ~new_n10136_;
  assign new_n6146_ = ~new_n10154_;
  assign new_n10147_ = new_n9595_ & new_n7376_;
  assign new_n6147_ = ~new_n10147_;
  assign new_n10288_ = D_REG_22_ | new_n10292_;
  assign new_n6148_ = ~new_n10288_;
  assign new_n10294_ = new_n10298_ | new_n10299_;
  assign new_n7065_ = ~new_n9244_;
  assign new_n7439_ = ~new_n10780_;
  assign new_n6149_ = ~new_n10294_;
  assign new_n10303_ = new_n10307_ | new_n10308_;
  assign new_n6150_ = ~new_n10303_;
  assign new_n10310_ = D_REG_25_ | new_n10314_;
  assign new_n6151_ = ~new_n10310_;
  assign new_n6152_ = ~new_n10336_;
  assign new_n10380_ = new_n7068_ | new_n6702_;
  assign new_n6153_ = ~new_n10380_;
  assign new_n10395_ = new_n7508_ & new_n10397_;
  assign new_n6154_ = ~new_n10395_;
  assign new_n7440_ = ~new_n10862_;
  assign new_n6155_ = ~new_n10406_;
  assign new_n10328_ = new_n6302_ | new_n6710_;
  assign new_n6156_ = ~new_n10328_;
  assign new_n6157_ = ~new_n10479_;
  assign new_n10480_ = new_n10338_ & new_n7521_;
  assign new_n6158_ = ~new_n10480_;
  assign new_n10484_ = new_n7067_ | new_n6712_;
  assign new_n6159_ = ~new_n10484_;
  assign new_n6160_ = ~new_n10493_;
  assign new_n6161_ = ~new_n10503_;
  assign new_n7441_ = ~new_n9912_;
  assign new_n6162_ = ~new_n10549_;
  assign new_n6163_ = ~new_n10551_;
  assign new_n6164_ = ~new_n10572_;
  assign new_n10580_ = new_n6305_ | new_n6715_;
  assign new_n6165_ = ~new_n10580_;
  assign new_n6166_ = ~new_n10626_;
  assign new_n6167_ = ~new_n10628_;
  assign new_n6168_ = ~new_n10630_;
  assign new_n10689_ = new_n7528_ | new_n9405_;
  assign new_n6169_ = ~new_n10689_;
  assign new_n7442_ = ~new_n8257_;
  assign new_n10325_ = new_n10698_ & B_REG;
  assign new_n6170_ = ~new_n10325_;
  assign new_n10705_ = DATAO_REG_31_ & new_n7566_;
  assign new_n6171_ = ~new_n10705_;
  assign new_n10715_ = DATAO_REG_30_ & new_n7566_;
  assign new_n6172_ = ~new_n10715_;
  assign new_n10721_ = DATAO_REG_29_ & new_n7566_;
  assign new_n6173_ = ~new_n10721_;
  assign new_n10731_ = DATAO_REG_28_ & new_n7566_;
  assign new_n6174_ = ~new_n10731_;
  assign new_n7443_ = ~new_n9290_;
  assign new_n10741_ = DATAO_REG_27_ & new_n7566_;
  assign new_n6175_ = ~new_n10741_;
  assign new_n10749_ = DATAO_REG_26_ & new_n7566_;
  assign new_n6176_ = ~new_n10749_;
  assign new_n10762_ = DATAO_REG_25_ & new_n7566_;
  assign new_n6177_ = ~new_n10762_;
  assign new_n10770_ = DATAO_REG_24_ & new_n7566_;
  assign new_n6178_ = ~new_n10770_;
  assign new_n10783_ = DATAO_REG_23_ & new_n7566_;
  assign new_n6179_ = ~new_n10783_;
  assign new_n9290_ = new_n9278_ & new_n9282_;
  assign new_n10791_ = DATAO_REG_22_ & new_n7566_;
  assign new_n6180_ = ~new_n10791_;
  assign new_n10802_ = DATAO_REG_21_ & new_n7566_;
  assign new_n6181_ = ~new_n10802_;
  assign new_n10811_ = DATAO_REG_20_ & new_n7566_;
  assign new_n6182_ = ~new_n10811_;
  assign new_n10823_ = DATAO_REG_19_ & new_n7566_;
  assign new_n6183_ = ~new_n10823_;
  assign new_n10831_ = DATAO_REG_18_ & new_n7566_;
  assign new_n6184_ = ~new_n10831_;
  assign new_n7444_ = ~new_n9265_;
  assign new_n10844_ = DATAO_REG_17_ & new_n7566_;
  assign new_n6185_ = ~new_n10844_;
  assign new_n10852_ = DATAO_REG_16_ & new_n7566_;
  assign new_n6186_ = ~new_n10852_;
  assign new_n10865_ = DATAO_REG_15_ & new_n7566_;
  assign new_n6187_ = ~new_n10865_;
  assign new_n10873_ = DATAO_REG_14_ & new_n7566_;
  assign new_n6188_ = ~new_n10873_;
  assign new_n10885_ = DATAO_REG_13_ & new_n7566_;
  assign new_n6189_ = ~new_n10885_;
  assign new_n7445_ = ~new_n8100_;
  assign new_n10893_ = DATAO_REG_12_ & new_n7566_;
  assign new_n6190_ = ~new_n10893_;
  assign new_n10906_ = DATAO_REG_11_ & new_n7566_;
  assign new_n6191_ = ~new_n10906_;
  assign new_n10914_ = DATAO_REG_10_ & new_n7566_;
  assign new_n6192_ = ~new_n10914_;
  assign new_n10927_ = DATAO_REG_9_ & new_n7566_;
  assign new_n6193_ = ~new_n10927_;
  assign new_n10935_ = DATAO_REG_8_ & new_n7566_;
  assign new_n6194_ = ~new_n10935_;
  assign new_n7446_ = ~new_n10596_;
  assign new_n10948_ = DATAO_REG_7_ & new_n7566_;
  assign new_n6195_ = ~new_n10948_;
  assign new_n10957_ = DATAO_REG_6_ & new_n7566_;
  assign new_n6196_ = ~new_n10957_;
  assign new_n10967_ = DATAO_REG_5_ & new_n7566_;
  assign new_n6197_ = ~new_n10967_;
  assign new_n10975_ = DATAO_REG_4_ & new_n7566_;
  assign new_n6198_ = ~new_n10975_;
  assign new_n10984_ = DATAO_REG_3_ & new_n7566_;
  assign new_n6199_ = ~new_n10984_;
  assign new_n7845_ = DATAI_26_ & new_n7551_;
  assign new_n10992_ = DATAO_REG_2_ & new_n7566_;
  assign new_n6200_ = ~new_n10992_;
  assign new_n11000_ = DATAO_REG_1_ & new_n7566_;
  assign new_n6201_ = ~new_n11000_;
  assign new_n11008_ = DATAO_REG_0_ & new_n7566_;
  assign new_n6202_ = ~new_n11008_;
  assign new_n11047_ = new_n7580_ & new_n11051_;
  assign new_n6203_ = ~new_n11047_;
  assign new_n11075_ = new_n6205_ & new_n11077_;
  assign new_n6204_ = ~new_n11075_;
  assign new_n7027_ = ~new_n8144_;
  assign new_n7066_ = ~new_n11117_;
  assign new_n7447_ = ~new_n7845_;
  assign new_n11076_ = new_n7586_ & new_n11080_;
  assign new_n6205_ = ~new_n11076_;
  assign new_n6206_ = ~new_n11095_;
  assign new_n11096_ = new_n11099_ & new_n7580_;
  assign new_n6207_ = ~new_n11096_;
  assign new_n11102_ = new_n11104_ & new_n11103_;
  assign new_n6208_ = ~new_n11102_;
  assign new_n11126_ = new_n9292_ | new_n9280_;
  assign new_n6209_ = ~new_n11126_;
  assign new_n11149_ = new_n7527_ | new_n9391_;
  assign new_n7448_ = ~new_n10649_;
  assign new_n6210_ = ~new_n11149_;
  assign new_n11169_ = new_n7586_ & new_n11173_;
  assign new_n6211_ = ~new_n11169_;
  assign new_n6212_ = ~new_n11189_;
  assign new_n11190_ = new_n11193_ & new_n7580_;
  assign new_n6213_ = ~new_n11190_;
  assign new_n11201_ = new_n7580_ & new_n11205_;
  assign new_n6214_ = ~new_n11201_;
  assign new_n11227_ = new_n6216_ & new_n11229_;
  assign new_n6215_ = ~new_n11227_;
  assign new_n7449_ = ~new_n10611_;
  assign new_n11228_ = new_n7586_ & new_n11232_;
  assign new_n6216_ = ~new_n11228_;
  assign new_n11239_ = new_n11243_ & new_n7580_;
  assign new_n6217_ = ~new_n11239_;
  assign new_n11265_ = new_n6219_ & new_n11267_;
  assign new_n6218_ = ~new_n11265_;
  assign new_n11266_ = new_n7586_ & new_n11270_;
  assign new_n6219_ = ~new_n11266_;
  assign new_n11277_ = new_n11281_ & new_n7580_;
  assign new_n6220_ = ~new_n11277_;
  assign new_n7450_ = ~new_n10119_;
  assign new_n6221_ = ~new_n11303_;
  assign new_n11340_ = new_n11341_ & new_n10596_;
  assign new_n6222_ = ~new_n11340_;
  assign new_n11308_ = new_n7580_ & new_n11346_;
  assign new_n6223_ = ~new_n11308_;
  assign new_n11349_ = new_n10652_ & new_n7495_;
  assign new_n6224_ = ~new_n11349_;
  assign new_n11361_ = new_n9464_ | new_n7467_;
  assign new_n6225_ = ~new_n11361_;
  assign new_n11378_ = new_n9536_ | new_n9484_;
  assign new_n9540_ = new_n11459_ & new_n10316_;
  assign new_n6226_ = ~new_n11378_;
  assign new_n11384_ = new_n7402_ & new_n7499_;
  assign new_n6227_ = ~new_n11384_;
  assign new_n11388_ = new_n9536_ | new_n7468_;
  assign new_n6228_ = ~new_n11388_;
  assign new_n11404_ = new_n9536_ | new_n7483_;
  assign new_n6229_ = ~new_n11404_;
  assign new_n11414_ = new_n9536_ | new_n9522_;
  assign new_n6230_ = ~new_n11414_;
  assign new_n11424_ = new_n9532_ | new_n9530_;
  assign new_n7451_ = ~new_n9540_;
  assign new_n6231_ = ~new_n11424_;
  assign new_n11445_ = new_n9376_ | new_n7466_;
  assign new_n6232_ = ~new_n11445_;
  assign new_n11450_ = new_n7481_ | new_n9338_;
  assign new_n6233_ = ~new_n11450_;
  assign new_n11454_ = new_n9329_ | new_n11447_;
  assign new_n6234_ = ~new_n11454_;
  assign new_n11468_ = new_n9361_ | new_n7465_;
  assign new_n6235_ = ~new_n11468_;
  assign new_n7802_ = new_n7519_ | new_n7559_;
  assign new_n7452_ = ~new_n10411_;
  assign new_n6236_ = ~new_n7802_;
  assign new_n6237_ = ~new_n7810_;
  assign new_n7822_ = new_n7457_ | new_n7559_;
  assign new_n6238_ = ~new_n7822_;
  assign new_n6239_ = ~new_n7829_;
  assign new_n7839_ = new_n7447_ | new_n7559_;
  assign new_n6240_ = ~new_n7839_;
  assign new_n6241_ = ~new_n7846_;
  assign new_n7856_ = new_n7512_ | new_n7559_;
  assign new_n6242_ = ~new_n7856_;
  assign new_n7453_ = ~new_n8968_;
  assign new_n6243_ = ~new_n7863_;
  assign new_n7873_ = new_n7454_ | new_n7559_;
  assign new_n6244_ = ~new_n7873_;
  assign new_n6245_ = ~new_n7880_;
  assign new_n7890_ = new_n7538_ | new_n7559_;
  assign new_n6246_ = ~new_n7890_;
  assign new_n6247_ = ~new_n7897_;
  assign new_n7907_ = new_n7395_ | new_n7559_;
  assign new_n6248_ = ~new_n7907_;
  assign new_n6249_ = ~new_n7914_;
  assign new_n7879_ = DATAI_24_ & new_n7551_;
  assign new_n7924_ = new_n7509_ | new_n7559_;
  assign new_n6250_ = ~new_n7924_;
  assign new_n6251_ = ~new_n7931_;
  assign new_n7941_ = new_n7385_ | new_n7559_;
  assign new_n6252_ = ~new_n7941_;
  assign new_n6253_ = ~new_n7948_;
  assign new_n7958_ = new_n7438_ | new_n7559_;
  assign new_n6254_ = ~new_n7958_;
  assign new_n6255_ = ~new_n7965_;
  assign new_n7975_ = new_n7456_ | new_n7559_;
  assign new_n7454_ = ~new_n7879_;
  assign new_n6256_ = ~new_n7975_;
  assign new_n6257_ = ~new_n7982_;
  assign new_n7992_ = new_n7536_ | new_n7559_;
  assign new_n6258_ = ~new_n7992_;
  assign new_n6259_ = ~new_n7999_;
  assign new_n8009_ = new_n7381_ | new_n7559_;
  assign new_n6260_ = ~new_n8009_;
  assign new_n6261_ = ~new_n8016_;
  assign new_n8026_ = new_n7532_ | new_n7559_;
  assign new_n6262_ = ~new_n8026_;
  assign new_n10478_ = new_n10527_ & new_n7110_;
  assign new_n7455_ = ~new_n7605_;
  assign new_n6263_ = ~new_n8033_;
  assign new_n8043_ = new_n7382_ | new_n7559_;
  assign new_n6264_ = ~new_n8043_;
  assign new_n6265_ = ~new_n8050_;
  assign new_n8060_ = new_n7437_ | new_n7559_;
  assign new_n6266_ = ~new_n8060_;
  assign new_n6267_ = ~new_n8067_;
  assign new_n8077_ = new_n7518_ | new_n7559_;
  assign new_n6268_ = ~new_n8077_;
  assign new_n6269_ = ~new_n8084_;
  assign new_n7456_ = ~new_n7981_;
  assign new_n8094_ = new_n7445_ | new_n7559_;
  assign new_n6270_ = ~new_n8094_;
  assign new_n6271_ = ~new_n8101_;
  assign new_n8111_ = new_n7380_ | new_n7559_;
  assign new_n6272_ = ~new_n8111_;
  assign new_n6273_ = ~new_n8120_;
  assign new_n8130_ = new_n7535_ | new_n7559_;
  assign new_n6274_ = ~new_n8130_;
  assign new_n6275_ = ~new_n8137_;
  assign new_n8147_ = new_n7393_ | new_n7559_;
  assign new_n7828_ = DATAI_27_ & new_n7551_;
  assign new_n6276_ = ~new_n8147_;
  assign new_n6277_ = ~new_n8155_;
  assign new_n8165_ = new_n7534_ | new_n7559_;
  assign new_n6278_ = ~new_n8165_;
  assign new_n6279_ = ~new_n8172_;
  assign new_n8182_ = new_n7379_ | new_n7559_;
  assign new_n6280_ = ~new_n8182_;
  assign new_n6281_ = ~new_n8190_;
  assign new_n8200_ = new_n7533_ | new_n7559_;
  assign new_n6282_ = ~new_n8200_;
  assign new_n7457_ = ~new_n7828_;
  assign new_n6283_ = ~new_n8207_;
  assign new_n6284_ = ~new_n8224_;
  assign new_n8233_ = new_n7531_ | new_n7559_;
  assign new_n6285_ = ~new_n8233_;
  assign new_n6286_ = ~new_n8240_;
  assign new_n8250_ = new_n7442_ | new_n7559_;
  assign new_n6287_ = ~new_n8250_;
  assign new_n6288_ = ~new_n8258_;
  assign new_n8268_ = new_n7549_ | new_n7559_;
  assign new_n6289_ = ~new_n8268_;
  assign new_n7458_ = ~new_n10375_;
  assign new_n6290_ = ~new_n8275_;
  assign new_n8437_ = new_n8439_ | new_n6701_;
  assign new_n6291_ = ~new_n8437_;
  assign new_n10430_ = new_n8584_ & new_n8564_;
  assign new_n6292_ = ~new_n10430_;
  assign new_n10434_ = new_n8710_ & new_n8685_;
  assign new_n6293_ = ~new_n10434_;
  assign new_n6294_ = ~new_n10426_;
  assign new_n10439_ = new_n10441_ & new_n7469_;
  assign new_n6295_ = ~new_n10439_;
  assign new_n7459_ = ~new_n10404_;
  assign new_n10443_ = new_n8467_ & new_n8439_;
  assign new_n6296_ = ~new_n10443_;
  assign new_n10450_ = new_n9089_ & new_n9057_;
  assign new_n6297_ = ~new_n10450_;
  assign new_n10453_ = new_n9208_ & new_n9185_;
  assign new_n6298_ = ~new_n10453_;
  assign new_n6299_ = ~new_n10446_;
  assign new_n10458_ = new_n10461_ & new_n8853_;
  assign new_n6300_ = ~new_n10458_;
  assign new_n10462_ = new_n8971_ & new_n8940_;
  assign new_n7460_ = ~new_n10652_;
  assign new_n6301_ = ~new_n10462_;
  assign new_n6302_ = ~new_n10466_;
  assign new_n6303_ = ~new_n10536_;
  assign new_n10582_ = new_n10590_ & new_n7525_;
  assign new_n6304_ = ~new_n10582_;
  assign new_n10599_ = new_n10604_ & new_n7135_;
  assign new_n6305_ = ~new_n10599_;
  assign new_n10620_ = new_n6307_ | new_n7098_;
  assign new_n6306_ = ~new_n10620_;
  assign new_n10632_ = new_n6308_ | new_n6717_;
  assign new_n7461_ = ~new_n8415_;
  assign new_n6307_ = ~new_n10632_;
  assign new_n6308_ = ~new_n10640_;
  assign new_n10655_ = new_n10668_ & new_n7485_;
  assign new_n6309_ = ~new_n10655_;
  assign new_n10681_ = new_n7479_ & new_n7515_;
  assign new_n6310_ = ~new_n10681_;
  assign new_n7588_ = new_n7580_ & new_n7189_;
  assign new_n6311_ = ~new_n7588_;
  assign new_n7602_ = new_n7580_ & new_n7190_;
  assign new_n6312_ = ~new_n7602_;
  assign new_n8415_ = DATAI_29_ & new_n7551_;
  assign new_n7627_ = new_n7580_ & new_n7191_;
  assign new_n6313_ = ~new_n7627_;
  assign new_n7641_ = new_n7642_ & new_n7586_;
  assign new_n6314_ = ~new_n7641_;
  assign new_n7670_ = new_n7671_ & new_n7586_;
  assign new_n6315_ = ~new_n7670_;
  assign new_n7685_ = new_n7686_ & new_n7586_;
  assign new_n6316_ = ~new_n7685_;
  assign new_n7740_ = new_n7741_ & new_n7586_;
  assign new_n6317_ = ~new_n7740_;
  assign new_n7462_ = ~new_n8472_;
  assign new_n8405_ = new_n7775_ & new_n8413_;
  assign new_n6318_ = ~new_n8405_;
  assign new_n6319_ = ~new_n8478_;
  assign new_n6320_ = ~new_n8498_;
  assign new_n8493_ = new_n7827_ & new_n8292_;
  assign new_n6321_ = ~new_n8493_;
  assign new_n6322_ = ~new_n8541_;
  assign new_n6323_ = ~new_n8591_;
  assign new_n6324_ = ~new_n8657_;
  assign new_n6325_ = ~new_n8719_;
  assign new_n7067_ = ~new_n10478_;
  assign new_n7463_ = ~new_n7617_;
  assign new_n8725_ = new_n8731_ & new_n7160_;
  assign new_n6326_ = ~new_n8725_;
  assign new_n8730_ = new_n7048_ & new_n7270_;
  assign new_n6327_ = ~new_n8730_;
  assign new_n6328_ = ~new_n8767_;
  assign new_n8798_ = new_n7101_ & new_n7333_;
  assign new_n6329_ = ~new_n8798_;
  assign new_n6330_ = ~new_n8830_;
  assign new_n8839_ = new_n7245_ & new_n7532_;
  assign new_n6331_ = ~new_n8839_;
  assign new_n7464_ = ~new_n7576_;
  assign new_n6332_ = ~new_n8885_;
  assign new_n6333_ = ~new_n8947_;
  assign new_n9099_ = new_n7097_ & new_n7334_;
  assign new_n6334_ = ~new_n9099_;
  assign new_n9164_ = new_n7102_ & new_n7033_;
  assign new_n6335_ = ~new_n9164_;
  assign new_n9562_ = new_n9567_ & new_n7290_;
  assign new_n6336_ = ~new_n9562_;
  assign new_n9566_ = new_n7050_ & new_n7412_;
  assign new_n6337_ = ~new_n9566_;
  assign new_n7465_ = ~new_n9359_;
  assign new_n9552_ = new_n8171_ & new_n7556_;
  assign new_n6338_ = ~new_n9552_;
  assign new_n9631_ = new_n7555_ & new_n8244_;
  assign new_n6339_ = ~new_n9631_;
  assign new_n9735_ = new_n7930_ & new_n7556_;
  assign new_n6340_ = ~new_n9735_;
  assign new_n9812_ = new_n7998_ & new_n7556_;
  assign new_n6341_ = ~new_n9812_;
  assign new_n9904_ = new_n9905_ & new_n7405_;
  assign new_n6342_ = ~new_n9904_;
  assign new_n7466_ = ~new_n9374_;
  assign new_n10031_ = new_n9740_ & new_n7071_;
  assign new_n6343_ = ~new_n10031_;
  assign new_n10107_ = new_n10122_ | new_n7444_;
  assign new_n6344_ = ~new_n10107_;
  assign new_n10108_ = new_n10122_ | new_n9265_;
  assign new_n6345_ = ~new_n10108_;
  assign new_n10115_ = new_n7256_ & new_n7547_;
  assign new_n6346_ = ~new_n10115_;
  assign new_n10183_ = new_n9640_ & new_n7074_;
  assign new_n6347_ = ~new_n10183_;
  assign new_n7467_ = ~new_n9462_;
  assign new_n10497_ = new_n8586_ & new_n7522_;
  assign new_n6348_ = ~new_n10497_;
  assign new_n10509_ = new_n10510_ & new_n7109_;
  assign new_n6349_ = ~new_n10509_;
  assign new_n10520_ = new_n9207_ & new_n7476_;
  assign new_n6350_ = ~new_n10520_;
  assign new_n6351_ = ~new_n10554_;
  assign new_n6352_ = ~new_n10558_;
  assign new_n10587_ = new_n7549_ & new_n10442_;
  assign new_n6353_ = ~new_n10587_;
  assign new_n7468_ = ~new_n9492_;
  assign new_n10699_ = new_n10704_ & new_n7547_;
  assign new_n6354_ = ~new_n10699_;
  assign new_n6355_ = ~new_n10757_;
  assign new_n6356_ = ~new_n10778_;
  assign new_n6357_ = ~new_n10819_;
  assign new_n6358_ = ~new_n10839_;
  assign new_n6359_ = ~new_n10860_;
  assign new_n6360_ = ~new_n10901_;
  assign new_n6361_ = ~new_n10922_;
  assign new_n6362_ = ~new_n10943_;
  assign new_n7469_ = ~new_n10337_;
  assign new_n11057_ = new_n11058_ & new_n7586_;
  assign new_n6363_ = ~new_n11057_;
  assign new_n11071_ = new_n11072_ & new_n7586_;
  assign new_n6364_ = ~new_n11071_;
  assign new_n11091_ = new_n11092_ & new_n7586_;
  assign new_n6365_ = ~new_n11091_;
  assign new_n11143_ = new_n7258_ & new_n7418_;
  assign new_n6366_ = ~new_n11143_;
  assign new_n11164_ = new_n11165_ & new_n7586_;
  assign new_n6367_ = ~new_n11164_;
  assign new_n7470_ = ~new_n8857_;
  assign new_n11185_ = new_n11186_ & new_n7586_;
  assign new_n6368_ = ~new_n11185_;
  assign new_n11211_ = new_n11212_ & new_n7586_;
  assign new_n6369_ = ~new_n11211_;
  assign new_n11223_ = new_n11224_ & new_n7586_;
  assign new_n6370_ = ~new_n11223_;
  assign new_n11249_ = new_n11250_ & new_n7586_;
  assign new_n6371_ = ~new_n11249_;
  assign new_n11261_ = new_n11262_ & new_n7586_;
  assign new_n6372_ = ~new_n11261_;
  assign new_n9061_ = new_n7534_ & new_n9075_;
  assign new_n11288_ = new_n11289_ & new_n7586_;
  assign new_n6373_ = ~new_n11288_;
  assign new_n11301_ = new_n11302_ & new_n7586_;
  assign new_n6374_ = ~new_n11301_;
  assign new_n11372_ = REG1_REG_7_ & new_n7146_;
  assign new_n6375_ = ~new_n11372_;
  assign new_n11396_ = IR_REG_5_ & new_n7276_;
  assign new_n6376_ = ~new_n11396_;
  assign new_n11408_ = REG1_REG_2_ & new_n7149_;
  assign new_n6377_ = ~new_n11408_;
  assign new_n7471_ = ~new_n9061_;
  assign new_n11435_ = new_n10119_ & new_n7551_;
  assign new_n6378_ = ~new_n11435_;
  assign new_n6379_ = ~new_n8425_;
  assign new_n6380_ = ~new_n8619_;
  assign new_n6381_ = ~new_n9283_;
  assign new_n6382_ = ~new_n10283_;
  assign new_n10519_ = new_n7508_ & new_n7472_;
  assign new_n6383_ = ~new_n10519_;
  assign new_n10605_ = new_n7473_ & new_n7475_;
  assign new_n6384_ = ~new_n10605_;
  assign new_n10384_ = new_n7281_ & new_n7399_;
  assign new_n7472_ = ~new_n10393_;
  assign new_n10634_ = new_n10342_ & new_n7413_;
  assign new_n6385_ = ~new_n10634_;
  assign new_n10637_ = new_n7477_ & new_n7422_;
  assign new_n6386_ = ~new_n10637_;
  assign new_n6387_ = ~new_n10733_;
  assign new_n6388_ = ~new_n10743_;
  assign new_n6389_ = ~new_n10751_;
  assign new_n6390_ = ~new_n10764_;
  assign new_n6391_ = ~new_n10772_;
  assign new_n6392_ = ~new_n10785_;
  assign new_n7473_ = ~new_n10396_;
  assign new_n6393_ = ~new_n10793_;
  assign new_n6394_ = ~new_n10804_;
  assign new_n6395_ = ~new_n10813_;
  assign new_n6396_ = ~new_n10825_;
  assign new_n6397_ = ~new_n10833_;
  assign new_n6398_ = ~new_n10846_;
  assign new_n6399_ = ~new_n10854_;
  assign new_n6400_ = ~new_n10867_;
  assign new_n6401_ = ~new_n10875_;
  assign new_n10881_ = REG3_REG_14_ | new_n10884_;
  assign new_n7474_ = ~new_n8615_;
  assign new_n6402_ = ~new_n10881_;
  assign new_n6403_ = ~new_n10887_;
  assign new_n6404_ = ~new_n10895_;
  assign new_n6405_ = ~new_n10908_;
  assign new_n6406_ = ~new_n10916_;
  assign new_n6407_ = ~new_n10929_;
  assign new_n6408_ = ~new_n10937_;
  assign new_n6409_ = ~new_n10950_;
  assign new_n6410_ = ~new_n10959_;
  assign new_n6411_ = ~new_n10969_;
  assign new_n9003_ = new_n7535_ & new_n9025_;
  assign new_n6412_ = ~new_n10977_;
  assign new_n6413_ = ~new_n10994_;
  assign new_n6414_ = ~new_n11002_;
  assign new_n6415_ = ~new_n11132_;
  assign new_n6416_ = ~new_n8426_;
  assign new_n6417_ = ~new_n8620_;
  assign new_n8672_ = new_n8665_ & new_n8750_;
  assign new_n6418_ = ~new_n8672_;
  assign new_n9191_ = new_n7369_ & new_n7531_;
  assign new_n6419_ = ~new_n9191_;
  assign new_n7475_ = ~new_n9003_;
  assign new_n9281_ = new_n7545_ & new_n7550_;
  assign new_n6420_ = ~new_n9281_;
  assign new_n9284_ = new_n10703_ & new_n7095_;
  assign new_n6421_ = ~new_n9284_;
  assign new_n6422_ = ~new_n10284_;
  assign new_n10606_ = new_n10525_ & new_n7520_;
  assign new_n6423_ = ~new_n10606_;
  assign new_n6424_ = ~new_n10638_;
  assign new_n6425_ = ~new_n10734_;
  assign new_n6426_ = ~new_n10744_;
  assign new_n10407_ = new_n7531_ & new_n8262_;
  assign new_n6427_ = ~new_n10752_;
  assign new_n6428_ = ~new_n10765_;
  assign new_n6429_ = ~new_n10773_;
  assign new_n6430_ = ~new_n10786_;
  assign new_n6431_ = ~new_n10794_;
  assign new_n6432_ = ~new_n10805_;
  assign new_n6433_ = ~new_n10814_;
  assign new_n6434_ = ~new_n10826_;
  assign new_n6435_ = ~new_n10834_;
  assign new_n6436_ = ~new_n10847_;
  assign new_n7476_ = ~new_n10407_;
  assign new_n6437_ = ~new_n10855_;
  assign new_n6438_ = ~new_n10868_;
  assign new_n6439_ = ~new_n10876_;
  assign new_n10883_ = REG3_REG_14_ & REG3_REG_13_;
  assign new_n6440_ = ~new_n10883_;
  assign new_n6441_ = ~new_n10888_;
  assign new_n6442_ = ~new_n10896_;
  assign new_n6443_ = ~new_n10909_;
  assign new_n6444_ = ~new_n10917_;
  assign new_n6445_ = ~new_n10930_;
  assign new_n8533_ = new_n8552_ & new_n7512_;
  assign new_n6446_ = ~new_n10938_;
  assign new_n6447_ = ~new_n10951_;
  assign new_n6448_ = ~new_n10960_;
  assign new_n6449_ = ~new_n10970_;
  assign new_n6450_ = ~new_n10978_;
  assign new_n6451_ = ~new_n10995_;
  assign new_n6452_ = ~new_n11003_;
  assign new_n6453_ = ~new_n11133_;
  assign new_n6454_ = ~new_n11385_;
  assign new_n6455_ = ~new_n11411_;
  assign new_n7477_ = ~new_n8533_;
  assign new_n6456_ = ~new_n11421_;
  assign new_n7736_ = new_n7121_ & new_n7737_;
  assign new_n6457_ = ~new_n7736_;
  assign new_n7789_ = REG2_REG_29_ & new_n7568_;
  assign new_n6458_ = ~new_n7789_;
  assign new_n7796_ = new_n7797_ & new_n7561_;
  assign new_n6459_ = ~new_n7796_;
  assign new_n8287_ = REG2_REG_0_ & new_n7568_;
  assign new_n6460_ = ~new_n8287_;
  assign new_n6461_ = ~new_n8297_;
  assign new_n7478_ = ~new_n10413_;
  assign new_n8465_ = new_n8466_ & new_n7560_;
  assign new_n6462_ = ~new_n8465_;
  assign new_n8477_ = new_n7806_ & new_n8413_;
  assign new_n6463_ = ~new_n8477_;
  assign new_n8507_ = new_n7826_ & new_n8413_;
  assign new_n6464_ = ~new_n8507_;
  assign new_n6465_ = ~new_n8519_;
  assign new_n8530_ = new_n8531_ & new_n7560_;
  assign new_n6466_ = ~new_n8530_;
  assign new_n8540_ = new_n7843_ & new_n8413_;
  assign new_n7068_ = ~new_n10384_;
  assign new_n7479_ = ~new_n10417_;
  assign new_n6467_ = ~new_n8540_;
  assign new_n8545_ = new_n8546_ & new_n8532_;
  assign new_n6468_ = ~new_n8545_;
  assign new_n8547_ = new_n8551_ & new_n7094_;
  assign new_n6469_ = ~new_n8547_;
  assign new_n8562_ = new_n8563_ & new_n7560_;
  assign new_n6470_ = ~new_n8562_;
  assign new_n8568_ = new_n7860_ & new_n8413_;
  assign new_n6471_ = ~new_n8568_;
  assign new_n8581_ = new_n8582_ & new_n7560_;
  assign new_n7480_ = ~new_n8429_;
  assign new_n6472_ = ~new_n8581_;
  assign new_n8590_ = new_n7877_ & new_n8413_;
  assign new_n6473_ = ~new_n8590_;
  assign new_n8607_ = new_n7560_ & new_n8608_;
  assign new_n6474_ = ~new_n8607_;
  assign new_n8633_ = new_n7894_ & new_n8413_;
  assign new_n6475_ = ~new_n8633_;
  assign new_n8648_ = new_n8649_ & new_n7560_;
  assign new_n6476_ = ~new_n8648_;
  assign new_n8656_ = new_n7911_ & new_n8413_;
  assign new_n7481_ = ~new_n9336_;
  assign new_n6477_ = ~new_n8656_;
  assign new_n8663_ = new_n8664_ & new_n8665_;
  assign new_n6478_ = ~new_n8663_;
  assign new_n8683_ = new_n8684_ & new_n7560_;
  assign new_n6479_ = ~new_n8683_;
  assign new_n8689_ = new_n7928_ & new_n8413_;
  assign new_n6480_ = ~new_n8689_;
  assign new_n8692_ = new_n8693_ & new_n7347_;
  assign new_n6481_ = ~new_n8692_;
  assign new_n8707_ = new_n8708_ & new_n7560_;
  assign new_n7482_ = ~new_n8628_;
  assign new_n6482_ = ~new_n8707_;
  assign new_n8718_ = new_n7945_ & new_n8413_;
  assign new_n6483_ = ~new_n8718_;
  assign new_n8723_ = new_n8724_ & new_n8710_;
  assign new_n6484_ = ~new_n8723_;
  assign new_n8740_ = new_n8741_ & new_n7560_;
  assign new_n6485_ = ~new_n8740_;
  assign new_n8746_ = new_n8413_ & new_n7962_;
  assign new_n6486_ = ~new_n8746_;
  assign new_n8759_ = new_n8760_ & new_n7560_;
  assign new_n7483_ = ~new_n9506_;
  assign new_n6487_ = ~new_n8759_;
  assign new_n8766_ = new_n7979_ & new_n8413_;
  assign new_n6488_ = ~new_n8766_;
  assign new_n8786_ = new_n8787_ & new_n7560_;
  assign new_n6489_ = ~new_n8786_;
  assign new_n8793_ = new_n8413_ & new_n7996_;
  assign new_n6490_ = ~new_n8793_;
  assign new_n8796_ = new_n8797_ & new_n8789_;
  assign new_n6491_ = ~new_n8796_;
  assign new_n8814_ = new_n8815_ & new_n7560_;
  assign new_n7484_ = ~new_n8713_;
  assign new_n6492_ = ~new_n8814_;
  assign new_n6493_ = ~new_n8817_;
  assign new_n8829_ = new_n8013_ & new_n8413_;
  assign new_n6494_ = ~new_n8829_;
  assign new_n8837_ = new_n8838_ & new_n8865_;
  assign new_n6495_ = ~new_n8837_;
  assign new_n8851_ = new_n8852_ & new_n7560_;
  assign new_n6496_ = ~new_n8851_;
  assign new_n8861_ = new_n8413_ & new_n8030_;
  assign new_n6497_ = ~new_n8861_;
  assign new_n10377_ = new_n7518_ & new_n8928_;
  assign new_n8878_ = new_n8879_ & new_n7560_;
  assign new_n6498_ = ~new_n8878_;
  assign new_n8884_ = new_n8047_ & new_n8413_;
  assign new_n6499_ = ~new_n8884_;
  assign new_n8897_ = new_n8898_ & new_n8100_;
  assign new_n6500_ = ~new_n8897_;
  assign new_n8908_ = new_n8909_ & new_n7560_;
  assign new_n6501_ = ~new_n8908_;
  assign new_n8915_ = new_n8413_ & new_n8064_;
  assign new_n6502_ = ~new_n8915_;
  assign new_n7485_ = ~new_n10377_;
  assign new_n8918_ = new_n8919_ & new_n8911_;
  assign new_n6503_ = ~new_n8918_;
  assign new_n6504_ = ~new_n8921_;
  assign new_n8937_ = new_n8938_ & new_n7560_;
  assign new_n6505_ = ~new_n8937_;
  assign new_n8946_ = new_n8081_ & new_n8413_;
  assign new_n6506_ = ~new_n8946_;
  assign new_n8961_ = new_n8962_ & new_n7560_;
  assign new_n6507_ = ~new_n8961_;
  assign new_n6508_ = ~new_n8964_;
  assign new_n7486_ = ~new_n8711_;
  assign new_n8976_ = new_n8413_ & new_n8098_;
  assign new_n6509_ = ~new_n8976_;
  assign new_n8987_ = new_n8988_ & new_n8154_;
  assign new_n6510_ = ~new_n8987_;
  assign new_n6511_ = ~new_n8998_;
  assign new_n9010_ = new_n9011_ & new_n8413_;
  assign new_n6512_ = ~new_n9010_;
  assign new_n9015_ = new_n9016_ & new_n9002_;
  assign new_n6513_ = ~new_n9015_;
  assign new_n6514_ = ~new_n9018_;
  assign new_n7487_ = ~new_n8535_;
  assign new_n9034_ = new_n9035_ & new_n7560_;
  assign new_n6515_ = ~new_n9034_;
  assign new_n9040_ = new_n8413_ & new_n8134_;
  assign new_n6516_ = ~new_n9040_;
  assign new_n9052_ = new_n9053_ & new_n7560_;
  assign new_n6517_ = ~new_n9052_;
  assign new_n6518_ = ~new_n9055_;
  assign new_n9067_ = new_n9068_ & new_n8413_;
  assign new_n6519_ = ~new_n9067_;
  assign new_n9087_ = new_n9088_ & new_n7560_;
  assign new_n9280_ = new_n9278_ & new_n7255_;
  assign new_n7586_ = new_n11345_ & new_n9265_;
  assign new_n6520_ = ~new_n9087_;
  assign new_n9095_ = new_n8413_ & new_n8169_;
  assign new_n6521_ = ~new_n9095_;
  assign new_n9097_ = new_n9098_ & new_n9089_;
  assign new_n6522_ = ~new_n9097_;
  assign new_n9115_ = new_n9116_ & new_n7560_;
  assign new_n6523_ = ~new_n9115_;
  assign new_n6524_ = ~new_n9118_;
  assign new_n9130_ = new_n9131_ & new_n8413_;
  assign new_n6525_ = ~new_n9130_;
  assign new_n7488_ = ~new_n7586_;
  assign new_n6526_ = ~new_n9139_;
  assign new_n6527_ = ~new_n9150_;
  assign new_n9160_ = new_n8413_ & new_n8204_;
  assign new_n6528_ = ~new_n9160_;
  assign new_n9162_ = new_n9163_ & new_n9154_;
  assign new_n6529_ = ~new_n9162_;
  assign new_n9182_ = new_n9183_ & new_n7560_;
  assign new_n6530_ = ~new_n9182_;
  assign new_n9189_ = new_n9190_ & new_n8413_;
  assign new_n6531_ = ~new_n9189_;
  assign new_n7489_ = ~new_n7664_;
  assign new_n9205_ = new_n9206_ & new_n7560_;
  assign new_n6532_ = ~new_n9205_;
  assign new_n9212_ = new_n8413_ & new_n8237_;
  assign new_n6533_ = ~new_n9212_;
  assign new_n9225_ = new_n9226_ & new_n7560_;
  assign new_n6534_ = ~new_n9225_;
  assign new_n9232_ = new_n9233_ & new_n8413_;
  assign new_n6535_ = ~new_n9232_;
  assign new_n9238_ = new_n9239_ & new_n9240_;
  assign new_n6536_ = ~new_n9238_;
  assign new_n7490_ = ~new_n7662_;
  assign new_n9253_ = new_n9254_ & new_n7560_;
  assign new_n6537_ = ~new_n9253_;
  assign new_n9260_ = new_n8413_ & new_n8272_;
  assign new_n6538_ = ~new_n9260_;
  assign new_n6539_ = ~new_n9267_;
  assign new_n6540_ = ~new_n9309_;
  assign new_n9318_ = new_n9319_ & new_n9313_;
  assign new_n6541_ = ~new_n9318_;
  assign new_n6542_ = ~new_n9325_;
  assign new_n6543_ = ~new_n9333_;
  assign new_n7491_ = ~new_n7683_;
  assign new_n9342_ = new_n9313_ & new_n7150_;
  assign new_n6544_ = ~new_n9342_;
  assign new_n6545_ = ~new_n9347_;
  assign new_n6546_ = ~new_n9356_;
  assign new_n9365_ = new_n9366_ & new_n9313_;
  assign new_n6547_ = ~new_n9365_;
  assign new_n6548_ = ~new_n9371_;
  assign new_n9380_ = new_n9381_ & new_n9313_;
  assign new_n6549_ = ~new_n9380_;
  assign new_n6550_ = ~new_n9386_;
  assign new_n7492_ = ~new_n7687_;
  assign new_n6551_ = ~new_n9395_;
  assign new_n6552_ = ~new_n9400_;
  assign new_n6553_ = ~new_n9409_;
  assign new_n6554_ = ~new_n9414_;
  assign new_n9423_ = new_n9424_ & new_n9313_;
  assign new_n6555_ = ~new_n9423_;
  assign new_n6556_ = ~new_n9429_;
  assign new_n9438_ = new_n9439_ & new_n9313_;
  assign new_n6557_ = ~new_n9438_;
  assign new_n6558_ = ~new_n9444_;
  assign new_n7493_ = ~new_n7643_;
  assign new_n9453_ = new_n9454_ & new_n9313_;
  assign new_n6559_ = ~new_n9453_;
  assign new_n6560_ = ~new_n9459_;
  assign new_n9468_ = new_n9469_ & new_n9313_;
  assign new_n6561_ = ~new_n9468_;
  assign new_n6562_ = ~new_n9474_;
  assign new_n9482_ = new_n9483_ & new_n9313_;
  assign new_n6563_ = ~new_n9482_;
  assign new_n6564_ = ~new_n9489_;
  assign new_n9498_ = new_n9313_ & new_n9499_;
  assign new_n7494_ = ~new_n11166_;
  assign new_n6565_ = ~new_n9498_;
  assign new_n6566_ = ~new_n9503_;
  assign new_n6567_ = ~new_n9512_;
  assign new_n9520_ = new_n9521_ & new_n9313_;
  assign new_n6568_ = ~new_n9520_;
  assign new_n6569_ = ~new_n9527_;
  assign new_n9578_ = new_n9579_ & new_n9554_;
  assign new_n6570_ = ~new_n9578_;
  assign new_n9592_ = new_n9593_ & new_n9554_;
  assign new_n6571_ = ~new_n9592_;
  assign new_n7495_ = ~new_n11282_;
  assign new_n9607_ = new_n9554_ & new_n9608_;
  assign new_n6572_ = ~new_n9607_;
  assign new_n9622_ = new_n9554_ & new_n9623_;
  assign new_n6573_ = ~new_n9622_;
  assign new_n9636_ = new_n9637_ & new_n9554_;
  assign new_n6574_ = ~new_n9636_;
  assign new_n9639_ = new_n9640_ & new_n7201_;
  assign new_n6575_ = ~new_n9639_;
  assign new_n9657_ = new_n9658_ & new_n9554_;
  assign new_n6576_ = ~new_n9657_;
  assign new_n7496_ = ~new_n11280_;
  assign new_n9672_ = new_n9673_ & new_n9554_;
  assign new_n6577_ = ~new_n9672_;
  assign new_n9697_ = new_n9681_ & new_n7828_;
  assign new_n6578_ = ~new_n9697_;
  assign new_n9707_ = new_n9708_ & new_n9554_;
  assign new_n6579_ = ~new_n9707_;
  assign new_n9720_ = new_n9721_ & new_n9554_;
  assign new_n6580_ = ~new_n9720_;
  assign new_n9758_ = new_n9554_ & new_n9759_;
  assign new_n6581_ = ~new_n9758_;
  assign new_n7069_ = ~new_n9280_;
  assign new_n7497_ = ~new_n11242_;
  assign new_n9772_ = new_n9773_ & new_n9554_;
  assign new_n6582_ = ~new_n9772_;
  assign new_n9786_ = new_n9554_ & new_n9787_;
  assign new_n6583_ = ~new_n9786_;
  assign new_n9800_ = new_n9554_ & new_n9801_;
  assign new_n6584_ = ~new_n9800_;
  assign new_n9833_ = new_n9554_ & new_n9834_;
  assign new_n6585_ = ~new_n9833_;
  assign new_n9848_ = new_n8222_ & new_n7555_;
  assign new_n6586_ = ~new_n9848_;
  assign new_n7498_ = ~new_n11204_;
  assign new_n9863_ = new_n9554_ & new_n9864_;
  assign new_n6587_ = ~new_n9863_;
  assign new_n9885_ = new_n9554_ & new_n9886_;
  assign new_n6588_ = ~new_n9885_;
  assign new_n9896_ = new_n9897_ & new_n9554_;
  assign new_n6589_ = ~new_n9896_;
  assign new_n6590_ = ~new_n9899_;
  assign new_n9922_ = new_n9923_ & new_n9554_;
  assign new_n6591_ = ~new_n9922_;
  assign new_n6592_ = ~new_n9937_;
  assign new_n7499_ = ~new_n11184_;
  assign new_n9942_ = new_n9943_ & new_n9944_;
  assign new_n6593_ = ~new_n9942_;
  assign new_n9956_ = new_n9957_ & new_n9554_;
  assign new_n6594_ = ~new_n9956_;
  assign new_n9967_ = new_n9968_ & new_n9554_;
  assign new_n6595_ = ~new_n9967_;
  assign new_n9982_ = new_n9554_ & new_n9983_;
  assign new_n6596_ = ~new_n9982_;
  assign new_n9996_ = new_n9997_ & new_n9554_;
  assign new_n6597_ = ~new_n9996_;
  assign new_n7500_ = ~new_n11263_;
  assign new_n9999_ = new_n9694_ & new_n7204_;
  assign new_n6598_ = ~new_n9999_;
  assign new_n10001_ = new_n7277_ & new_n7345_;
  assign new_n6599_ = ~new_n10001_;
  assign new_n10040_ = new_n9745_ & new_n7278_;
  assign new_n6600_ = ~new_n10040_;
  assign new_n10048_ = new_n9681_ & new_n7964_;
  assign new_n6601_ = ~new_n10048_;
  assign new_n6602_ = ~new_n10050_;
  assign new_n10061_ = new_n9821_ & new_n7273_;
  assign new_n7501_ = ~new_n11225_;
  assign new_n6603_ = ~new_n10061_;
  assign new_n10125_ = new_n10126_ & new_n9554_;
  assign new_n6604_ = ~new_n10125_;
  assign new_n6605_ = ~new_n10132_;
  assign new_n10169_ = new_n7157_ & new_n7227_;
  assign new_n6606_ = ~new_n10169_;
  assign new_n10176_ = new_n10177_ & new_n9986_;
  assign new_n6607_ = ~new_n10176_;
  assign new_n10182_ = new_n9681_ & new_n9172_;
  assign new_n6608_ = ~new_n10182_;
  assign new_n7502_ = ~new_n11187_;
  assign new_n10192_ = new_n7279_ & new_n7346_;
  assign new_n6609_ = ~new_n10192_;
  assign new_n10321_ = new_n10323_ & new_n8432_;
  assign new_n6610_ = ~new_n10321_;
  assign new_n10331_ = new_n10332_ & new_n8450_;
  assign new_n6611_ = ~new_n10331_;
  assign new_n6612_ = ~new_n10333_;
  assign new_n6613_ = ~new_n10391_;
  assign new_n10514_ = new_n10515_ & new_n10516_;
  assign new_n6614_ = ~new_n10514_;
  assign new_n7503_ = ~new_n11093_;
  assign new_n10518_ = new_n7197_ & new_n10390_;
  assign new_n6615_ = ~new_n10518_;
  assign new_n6616_ = ~new_n10523_;
  assign new_n10636_ = new_n10352_ & new_n8615_;
  assign new_n6617_ = ~new_n10636_;
  assign new_n10666_ = new_n9419_ & new_n9536_;
  assign new_n6618_ = ~new_n10666_;
  assign new_n10688_ = new_n9405_ & new_n9536_;
  assign new_n6619_ = ~new_n10688_;
  assign new_n10696_ = new_n9434_ & new_n9536_;
  assign new_n7504_ = ~new_n11073_;
  assign new_n6620_ = ~new_n10696_;
  assign new_n10711_ = REG0_REG_31_ & new_n7562_;
  assign new_n6621_ = ~new_n10711_;
  assign new_n10720_ = REG0_REG_30_ & new_n7562_;
  assign new_n6622_ = ~new_n10720_;
  assign new_n11031_ = new_n7586_ & new_n11032_;
  assign new_n6623_ = ~new_n11031_;
  assign new_n11108_ = new_n11106_ & IR_REG_0_;
  assign new_n6624_ = ~new_n11108_;
  assign new_n11113_ = new_n9681_ & new_n9235_;
  assign new_n7505_ = ~new_n7767_;
  assign new_n6625_ = ~new_n11113_;
  assign new_n11119_ = new_n9282_ & new_n11129_;
  assign new_n6626_ = ~new_n11119_;
  assign new_n11123_ = new_n9235_ & new_n7557_;
  assign new_n6627_ = ~new_n11123_;
  assign new_n11148_ = new_n9391_ & new_n9536_;
  assign new_n6628_ = ~new_n11148_;
  assign new_n11306_ = new_n9449_ & new_n9536_;
  assign new_n6629_ = ~new_n11306_;
  assign new_n11360_ = new_n9464_ & new_n9536_;
  assign new_n7506_ = ~new_n9255_;
  assign new_n6630_ = ~new_n11360_;
  assign new_n11363_ = new_n7144_ & new_n11364_;
  assign new_n6631_ = ~new_n11363_;
  assign new_n11377_ = new_n9536_ & new_n9478_;
  assign new_n6632_ = ~new_n11377_;
  assign new_n11399_ = new_n7147_ & new_n11400_;
  assign new_n6633_ = ~new_n11399_;
  assign new_n11403_ = new_n9536_ & new_n9508_;
  assign new_n6634_ = ~new_n11403_;
  assign new_n11437_ = new_n7551_ & new_n7443_;
  assign new_n8515_ = new_n7239_ & new_n7447_;
  assign new_n7507_ = ~new_n8255_;
  assign new_n6635_ = ~new_n11437_;
  assign new_n11444_ = new_n9376_ & new_n9536_;
  assign new_n6636_ = ~new_n11444_;
  assign new_n11449_ = new_n9338_ & new_n9536_;
  assign new_n6637_ = ~new_n11449_;
  assign new_n11453_ = new_n9329_ & new_n9536_;
  assign new_n6638_ = ~new_n11453_;
  assign new_n11463_ = new_n9351_ & new_n9536_;
  assign new_n6639_ = ~new_n11463_;
  assign new_n11467_ = new_n9361_ & new_n9536_;
  assign new_n7508_ = ~new_n9122_;
  assign new_n6640_ = ~new_n11467_;
  assign new_n6641_ = ~new_n7803_;
  assign new_n6642_ = ~new_n7811_;
  assign new_n6643_ = ~new_n7823_;
  assign new_n6644_ = ~new_n7830_;
  assign new_n6645_ = ~new_n7840_;
  assign new_n6646_ = ~new_n7847_;
  assign new_n6647_ = ~new_n7857_;
  assign new_n6648_ = ~new_n7864_;
  assign new_n6649_ = ~new_n7874_;
  assign new_n7930_ = DATAI_21_ & new_n7551_;
  assign new_n6650_ = ~new_n7881_;
  assign new_n6651_ = ~new_n7891_;
  assign new_n6652_ = ~new_n7898_;
  assign new_n6653_ = ~new_n7908_;
  assign new_n6654_ = ~new_n7915_;
  assign new_n6655_ = ~new_n7925_;
  assign new_n6656_ = ~new_n7932_;
  assign new_n6657_ = ~new_n7942_;
  assign new_n6658_ = ~new_n7949_;
  assign new_n6659_ = ~new_n7959_;
  assign new_n7509_ = ~new_n7930_;
  assign new_n6660_ = ~new_n7966_;
  assign new_n6661_ = ~new_n7976_;
  assign new_n6662_ = ~new_n7983_;
  assign new_n6663_ = ~new_n7993_;
  assign new_n6664_ = ~new_n8000_;
  assign new_n6665_ = ~new_n8010_;
  assign new_n6666_ = ~new_n8017_;
  assign new_n6667_ = ~new_n8027_;
  assign new_n6668_ = ~new_n8034_;
  assign new_n6669_ = ~new_n8044_;
  assign new_n7510_ = ~new_n7739_;
  assign new_n6670_ = ~new_n8051_;
  assign new_n6671_ = ~new_n8061_;
  assign new_n6672_ = ~new_n8068_;
  assign new_n6673_ = ~new_n8078_;
  assign new_n6674_ = ~new_n8085_;
  assign new_n6675_ = ~new_n8095_;
  assign new_n6676_ = ~new_n8102_;
  assign new_n6677_ = ~new_n8112_;
  assign new_n6678_ = ~new_n8121_;
  assign new_n6679_ = ~new_n8131_;
  assign new_n7511_ = ~new_n10593_;
  assign new_n6680_ = ~new_n8138_;
  assign new_n6681_ = ~new_n8148_;
  assign new_n6682_ = ~new_n8156_;
  assign new_n6683_ = ~new_n8166_;
  assign new_n6684_ = ~new_n8173_;
  assign new_n6685_ = ~new_n8183_;
  assign new_n6686_ = ~new_n8191_;
  assign new_n6687_ = ~new_n8201_;
  assign new_n6688_ = ~new_n8208_;
  assign new_n6689_ = ~new_n8218_;
  assign new_n7862_ = DATAI_25_ & new_n7551_;
  assign new_n6690_ = ~new_n8225_;
  assign new_n6691_ = ~new_n8234_;
  assign new_n6692_ = ~new_n8241_;
  assign new_n6693_ = ~new_n8251_;
  assign new_n6694_ = ~new_n8259_;
  assign new_n6695_ = ~new_n8269_;
  assign new_n6696_ = ~new_n8276_;
  assign new_n8412_ = new_n7265_ | new_n6698_;
  assign new_n6697_ = ~new_n8412_;
  assign new_n6698_ = ~new_n7781_;
  assign new_n7512_ = ~new_n7862_;
  assign new_n8438_ = new_n7352_ | new_n6700_;
  assign new_n6699_ = ~new_n8438_;
  assign new_n6700_ = ~new_n8440_;
  assign new_n6701_ = ~new_n8445_;
  assign new_n6702_ = ~new_n10385_;
  assign new_n6703_ = ~new_n10427_;
  assign new_n10431_ = new_n8650_ & new_n8614_;
  assign new_n6704_ = ~new_n10431_;
  assign new_n10435_ = new_n8762_ & new_n8742_;
  assign new_n6705_ = ~new_n10435_;
  assign new_n7513_ = ~new_n7646_;
  assign new_n10444_ = new_n8532_ & new_n8503_;
  assign new_n6706_ = ~new_n10444_;
  assign new_n6707_ = ~new_n10447_;
  assign new_n10451_ = new_n9154_ & new_n9120_;
  assign new_n6708_ = ~new_n10451_;
  assign new_n10459_ = new_n8911_ & new_n8880_;
  assign new_n6709_ = ~new_n10459_;
  assign new_n6710_ = ~new_n10467_;
  assign new_n10486_ = new_n7543_ & new_n7539_;
  assign new_n6711_ = ~new_n10486_;
  assign new_n7514_ = ~new_n8502_;
  assign new_n6712_ = ~new_n10487_;
  assign new_n10537_ = new_n10538_ & new_n10539_;
  assign new_n6713_ = ~new_n10537_;
  assign new_n6714_ = ~new_n10583_;
  assign new_n10600_ = new_n10601_ & new_n10542_;
  assign new_n6715_ = ~new_n10600_;
  assign new_n6716_ = ~new_n10621_;
  assign new_n6717_ = ~new_n10641_;
  assign new_n6718_ = ~new_n10504_;
  assign new_n10682_ = new_n10361_ & new_n7546_;
  assign new_n7070_ = ~new_n8515_;
  assign new_n7515_ = ~new_n8854_;
  assign new_n6719_ = ~new_n10682_;
  assign new_n6720_ = ~new_n7571_;
  assign new_n6721_ = ~new_n7593_;
  assign new_n6722_ = ~new_n7612_;
  assign new_n6723_ = ~new_n7631_;
  assign new_n6724_ = ~new_n7652_;
  assign new_n6725_ = ~new_n7674_;
  assign new_n6726_ = ~new_n7696_;
  assign new_n6727_ = ~new_n7769_;
  assign new_n6728_ = ~new_n7777_;
  assign new_n7516_ = ~new_n10617_;
  assign new_n6729_ = ~new_n7785_;
  assign new_n6730_ = ~new_n9011_;
  assign new_n6731_ = ~new_n9068_;
  assign new_n6732_ = ~new_n9131_;
  assign new_n6733_ = ~new_n9190_;
  assign new_n6734_ = ~new_n9233_;
  assign new_n6735_ = ~new_n8283_;
  assign new_n8288_ = new_n8289_ & new_n7411_;
  assign new_n6736_ = ~new_n8288_;
  assign new_n6737_ = ~new_n8423_;
  assign new_n7517_ = ~new_n10614_;
  assign new_n6738_ = ~new_n8460_;
  assign new_n6739_ = ~new_n8489_;
  assign new_n6740_ = ~new_n8496_;
  assign new_n6741_ = ~new_n8525_;
  assign new_n6742_ = ~new_n8549_;
  assign new_n6743_ = ~new_n8557_;
  assign new_n6744_ = ~new_n8576_;
  assign new_n6745_ = ~new_n8602_;
  assign new_n6746_ = ~new_n8610_;
  assign new_n6747_ = ~new_n8643_;
  assign new_n7518_ = ~new_n8083_;
  assign new_n6748_ = ~new_n8678_;
  assign new_n6749_ = ~new_n8702_;
  assign new_n6750_ = ~new_n8735_;
  assign new_n6751_ = ~new_n8754_;
  assign new_n6752_ = ~new_n8781_;
  assign new_n6753_ = ~new_n8801_;
  assign new_n6754_ = ~new_n8809_;
  assign new_n6755_ = ~new_n8846_;
  assign new_n6756_ = ~new_n8873_;
  assign new_n6757_ = ~new_n8903_;
  assign new_n7519_ = ~new_n7808_;
  assign new_n6758_ = ~new_n8924_;
  assign new_n6759_ = ~new_n8932_;
  assign new_n6760_ = ~new_n8956_;
  assign new_n6761_ = ~new_n8993_;
  assign new_n6762_ = ~new_n9021_;
  assign new_n6763_ = ~new_n9029_;
  assign new_n6764_ = ~new_n9047_;
  assign new_n6765_ = ~new_n9082_;
  assign new_n6766_ = ~new_n9102_;
  assign new_n6767_ = ~new_n9110_;
  assign new_n7808_ = DATAI_28_ & new_n7551_;
  assign new_n6768_ = ~new_n9145_;
  assign new_n6769_ = ~new_n9167_;
  assign new_n6770_ = ~new_n9177_;
  assign new_n6771_ = ~new_n9200_;
  assign new_n6772_ = ~new_n9220_;
  assign new_n6773_ = ~new_n9248_;
  assign new_n6774_ = ~new_n9275_;
  assign new_n9279_ = new_n11129_ & new_n7545_;
  assign new_n6775_ = ~new_n9279_;
  assign new_n9304_ = new_n9313_ & new_n9305_;
  assign new_n9125_ = new_n7533_ & new_n9173_;
  assign new_n6776_ = ~new_n9304_;
  assign new_n9539_ = new_n7443_ & new_n7451_;
  assign new_n6777_ = ~new_n9539_;
  assign new_n9542_ = new_n9543_ & new_n7138_;
  assign new_n6778_ = ~new_n9542_;
  assign new_n6779_ = ~new_n9555_;
  assign new_n6780_ = ~new_n9570_;
  assign new_n9585_ = new_n9586_ & new_n7127_;
  assign new_n6781_ = ~new_n9585_;
  assign new_n6782_ = ~new_n9599_;
  assign new_n7520_ = ~new_n9125_;
  assign new_n9614_ = new_n9615_ & new_n7141_;
  assign new_n6783_ = ~new_n9614_;
  assign new_n6784_ = ~new_n9628_;
  assign new_n6785_ = ~new_n9642_;
  assign new_n9650_ = new_n9651_ & new_n7128_;
  assign new_n6786_ = ~new_n9650_;
  assign new_n6787_ = ~new_n9664_;
  assign new_n9699_ = new_n9700_ & new_n7139_;
  assign new_n6788_ = ~new_n9699_;
  assign new_n6789_ = ~new_n9714_;
  assign new_n7521_ = ~new_n8419_;
  assign new_n6790_ = ~new_n9728_;
  assign new_n6791_ = ~new_n9737_;
  assign new_n6792_ = ~new_n9742_;
  assign new_n9750_ = new_n9751_ & new_n7143_;
  assign new_n6793_ = ~new_n9750_;
  assign new_n6794_ = ~new_n9764_;
  assign new_n9779_ = new_n9780_ & new_n7129_;
  assign new_n6795_ = ~new_n9779_;
  assign new_n9792_ = new_n9793_ & new_n7136_;
  assign new_n6796_ = ~new_n9792_;
  assign new_n7522_ = ~new_n10433_;
  assign new_n9806_ = new_n9807_ & new_n7130_;
  assign new_n6797_ = ~new_n9806_;
  assign new_n6798_ = ~new_n9814_;
  assign new_n6799_ = ~new_n9819_;
  assign new_n6800_ = ~new_n9825_;
  assign new_n9840_ = new_n9841_ & new_n7111_;
  assign new_n6801_ = ~new_n9840_;
  assign new_n9855_ = new_n9856_ & new_n7140_;
  assign new_n6802_ = ~new_n9855_;
  assign new_n6803_ = ~new_n9870_;
  assign new_n7071_ = ~new_n9747_;
  assign new_n10412_ = new_n7536_ & new_n8774_;
  assign new_n6804_ = ~new_n9877_;
  assign new_n9889_ = new_n9890_ & new_n7131_;
  assign new_n6805_ = ~new_n9889_;
  assign new_n6806_ = ~new_n9907_;
  assign new_n6807_ = ~new_n9914_;
  assign new_n9929_ = new_n9930_ & new_n7142_;
  assign new_n6808_ = ~new_n9929_;
  assign new_n6809_ = ~new_n9950_;
  assign new_n9960_ = new_n9961_ & new_n7132_;
  assign new_n6810_ = ~new_n9960_;
  assign new_n7523_ = ~new_n10412_;
  assign new_n9974_ = new_n9975_ & new_n7137_;
  assign new_n6811_ = ~new_n9974_;
  assign new_n6812_ = ~new_n9988_;
  assign new_n6813_ = ~new_n10002_;
  assign new_n10103_ = new_n10104_ & new_n7133_;
  assign new_n6814_ = ~new_n10103_;
  assign new_n6815_ = ~new_n10118_;
  assign new_n6816_ = ~new_n10372_;
  assign new_n6817_ = ~new_n10399_;
  assign new_n10403_ = new_n7459_ & new_n10405_;
  assign new_n7524_ = ~new_n8443_;
  assign new_n6818_ = ~new_n10403_;
  assign new_n6819_ = ~new_n10472_;
  assign new_n10507_ = new_n7541_ & new_n7356_;
  assign new_n6820_ = ~new_n10507_;
  assign new_n10541_ = new_n10578_ & new_n10542_;
  assign new_n6821_ = ~new_n10541_;
  assign new_n10562_ = new_n10578_ & new_n10563_;
  assign new_n6822_ = ~new_n10562_;
  assign new_n6823_ = ~new_n10565_;
  assign new_n6824_ = ~new_n10569_;
  assign new_n7525_ = ~new_n9155_;
  assign new_n10701_ = new_n9265_ & new_n11106_;
  assign new_n6825_ = ~new_n10701_;
  assign new_n6826_ = ~new_n10724_;
  assign new_n6827_ = ~new_n10987_;
  assign new_n6828_ = ~new_n11011_;
  assign new_n11020_ = new_n11021_ & new_n7432_;
  assign new_n6829_ = ~new_n11020_;
  assign new_n11023_ = REG2_REG_0_ & new_n9530_;
  assign new_n6830_ = ~new_n11023_;
  assign new_n6831_ = ~new_n11025_;
  assign new_n7526_ = ~new_n8623_;
  assign new_n6832_ = ~new_n11041_;
  assign new_n6833_ = ~new_n11062_;
  assign new_n11082_ = new_n11083_ & new_n7111_;
  assign new_n6834_ = ~new_n11082_;
  assign new_n6835_ = ~new_n11155_;
  assign new_n6836_ = ~new_n11175_;
  assign new_n6837_ = ~new_n11196_;
  assign new_n6838_ = ~new_n11215_;
  assign new_n6839_ = ~new_n11234_;
  assign new_n6840_ = ~new_n11253_;
  assign new_n7527_ = ~new_n9389_;
  assign new_n6841_ = ~new_n11272_;
  assign new_n6842_ = ~new_n11292_;
  assign new_n6843_ = ~new_n11379_;
  assign new_n6844_ = ~new_n11415_;
  assign new_n6845_ = ~new_n7570_;
  assign new_n6846_ = ~new_n7592_;
  assign new_n6847_ = ~new_n7611_;
  assign new_n6848_ = ~new_n7630_;
  assign new_n6849_ = ~new_n7651_;
  assign new_n6850_ = ~new_n7673_;
  assign new_n7528_ = ~new_n9403_;
  assign new_n6851_ = ~new_n7695_;
  assign new_n6852_ = ~new_n7768_;
  assign new_n6853_ = ~new_n7776_;
  assign new_n6854_ = ~new_n7784_;
  assign new_n6855_ = ~new_n8282_;
  assign new_n6856_ = ~new_n8422_;
  assign new_n6857_ = ~new_n8459_;
  assign new_n6858_ = ~new_n8495_;
  assign new_n6859_ = ~new_n8488_;
  assign new_n6860_ = ~new_n8524_;
  assign new_n7529_ = ~new_n10376_;
  assign new_n6861_ = ~new_n8556_;
  assign new_n6862_ = ~new_n8575_;
  assign new_n6863_ = ~new_n8609_;
  assign new_n6864_ = ~new_n8601_;
  assign new_n6865_ = ~new_n8642_;
  assign new_n6866_ = ~new_n8670_;
  assign new_n6867_ = ~new_n8677_;
  assign new_n6868_ = ~new_n8701_;
  assign new_n6869_ = ~new_n8734_;
  assign new_n6870_ = ~new_n8753_;
  assign new_n7530_ = ~new_n8618_;
  assign new_n6871_ = ~new_n8780_;
  assign new_n6872_ = ~new_n8808_;
  assign new_n6873_ = ~new_n8845_;
  assign new_n6874_ = ~new_n8872_;
  assign new_n6875_ = ~new_n8902_;
  assign new_n6876_ = ~new_n8931_;
  assign new_n6877_ = ~new_n8955_;
  assign new_n6878_ = ~new_n8992_;
  assign new_n6879_ = ~new_n9028_;
  assign new_n6880_ = ~new_n9046_;
  assign new_n7531_ = ~new_n8239_;
  assign new_n6881_ = ~new_n9081_;
  assign new_n6882_ = ~new_n9109_;
  assign new_n6883_ = ~new_n9144_;
  assign new_n6884_ = ~new_n9176_;
  assign new_n6885_ = ~new_n9199_;
  assign new_n6886_ = ~new_n9219_;
  assign new_n6887_ = ~new_n9247_;
  assign new_n6888_ = ~new_n9274_;
  assign new_n6889_ = ~new_n9541_;
  assign new_n6890_ = ~new_n9569_;
  assign new_n7028_ = ~new_n8162_;
  assign new_n7072_ = ~new_n9822_;
  assign new_n7532_ = ~new_n8032_;
  assign new_n6891_ = ~new_n9584_;
  assign new_n6892_ = ~new_n9598_;
  assign new_n6893_ = ~new_n9613_;
  assign new_n6894_ = ~new_n9627_;
  assign new_n6895_ = ~new_n9649_;
  assign new_n6896_ = ~new_n9663_;
  assign new_n6897_ = ~new_n9698_;
  assign new_n6898_ = ~new_n9713_;
  assign new_n6899_ = ~new_n9727_;
  assign new_n6900_ = ~new_n9749_;
  assign new_n7533_ = ~new_n8206_;
  assign new_n6901_ = ~new_n9763_;
  assign new_n6902_ = ~new_n9778_;
  assign new_n6903_ = ~new_n9791_;
  assign new_n6904_ = ~new_n9805_;
  assign new_n6905_ = ~new_n9824_;
  assign new_n6906_ = ~new_n9839_;
  assign new_n6907_ = ~new_n9854_;
  assign new_n6908_ = ~new_n9869_;
  assign new_n6909_ = ~new_n9876_;
  assign new_n6910_ = ~new_n9888_;
  assign new_n7534_ = ~new_n8171_;
  assign new_n9906_ = new_n7405_ & new_n7274_;
  assign new_n6911_ = ~new_n9906_;
  assign new_n6912_ = ~new_n9913_;
  assign new_n6913_ = ~new_n9928_;
  assign new_n6914_ = ~new_n9949_;
  assign new_n6915_ = ~new_n9959_;
  assign new_n6916_ = ~new_n9973_;
  assign new_n6917_ = ~new_n9987_;
  assign new_n6918_ = ~new_n10102_;
  assign new_n10117_ = new_n7159_ & new_n7451_;
  assign new_n7535_ = ~new_n8136_;
  assign new_n6919_ = ~new_n10117_;
  assign new_n10282_ = new_n7159_ & new_n7386_;
  assign new_n6920_ = ~new_n10282_;
  assign new_n6921_ = ~new_n10371_;
  assign new_n10398_ = new_n7525_ & new_n7520_;
  assign new_n6922_ = ~new_n10398_;
  assign new_n6923_ = ~new_n10471_;
  assign new_n10506_ = new_n7452_ & new_n7470_;
  assign new_n6924_ = ~new_n10506_;
  assign new_n6925_ = ~new_n10540_;
  assign new_n7536_ = ~new_n7998_;
  assign new_n10568_ = new_n7478_ & new_n7523_;
  assign new_n6926_ = ~new_n10568_;
  assign new_n6927_ = ~new_n10564_;
  assign new_n10561_ = new_n7546_ & new_n7479_;
  assign new_n6928_ = ~new_n10561_;
  assign new_n6929_ = ~new_n10723_;
  assign new_n6930_ = ~new_n10986_;
  assign new_n11010_ = new_n11014_ & new_n11015_;
  assign new_n6931_ = ~new_n11010_;
  assign new_n11024_ = new_n11028_ & new_n11029_;
  assign new_n7537_ = ~new_n7689_;
  assign new_n6932_ = ~new_n11024_;
  assign new_n6933_ = ~new_n11040_;
  assign new_n6934_ = ~new_n11061_;
  assign new_n6935_ = ~new_n11081_;
  assign new_n6936_ = ~new_n11154_;
  assign new_n6937_ = ~new_n11174_;
  assign new_n6938_ = ~new_n11195_;
  assign new_n6939_ = ~new_n11214_;
  assign new_n6940_ = ~new_n11233_;
  assign new_n6941_ = ~new_n11252_;
  assign new_n7538_ = ~new_n7896_;
  assign new_n6942_ = ~new_n11271_;
  assign new_n6943_ = ~new_n11291_;
  assign new_n6944_ = ~new_n8451_;
  assign new_n6945_ = ~new_n8863_;
  assign new_n8888_ = new_n7156_ & new_n7022_;
  assign new_n6946_ = ~new_n8888_;
  assign new_n6947_ = ~new_n9684_;
  assign new_n9709_ = new_n7157_ & new_n7161_;
  assign new_n6948_ = ~new_n9709_;
  assign new_n9722_ = new_n7134_ & new_n7075_;
  assign new_n7896_ = DATAI_23_ & new_n7551_;
  assign new_n6949_ = ~new_n9722_;
  assign new_n9774_ = new_n7299_ & new_n7277_;
  assign new_n6950_ = ~new_n9774_;
  assign new_n9958_ = new_n7301_ & new_n7279_;
  assign new_n6951_ = ~new_n9958_;
  assign new_n6952_ = ~new_n10423_;
  assign new_n10739_ = REG3_REG_27_ & new_n10740_;
  assign new_n6953_ = ~new_n10739_;
  assign new_n10965_ = REG3_REG_5_ & new_n10966_;
  assign new_n6954_ = ~new_n10965_;
  assign new_n7539_ = ~new_n8442_;
  assign new_n6955_ = ~new_n8709_;
  assign new_n8939_ = new_n7198_ & new_n7109_;
  assign new_n6956_ = ~new_n8939_;
  assign new_n6957_ = ~new_n9676_;
  assign new_n6958_ = ~new_n9689_;
  assign new_n6959_ = ~new_n10015_;
  assign new_n6960_ = ~new_n10023_;
  assign new_n6961_ = ~new_n10076_;
  assign new_n6962_ = ~new_n10081_;
  assign new_n6963_ = ~new_n10091_;
  assign new_n7540_ = ~new_n7657_;
  assign new_n6964_ = ~new_n10140_;
  assign new_n6965_ = ~new_n10215_;
  assign new_n6966_ = ~new_n10221_;
  assign new_n6967_ = ~new_n10248_;
  assign new_n6968_ = ~new_n10260_;
  assign new_n6969_ = ~new_n10271_;
  assign new_n6970_ = ~new_n11115_;
  assign new_n9624_ = new_n7271_ & new_n7291_;
  assign new_n6971_ = ~new_n9624_;
  assign new_n9760_ = new_n7405_ & new_n7416_;
  assign new_n7073_ = ~new_n9695_;
  assign new_n7541_ = ~new_n8821_;
  assign new_n6972_ = ~new_n9760_;
  assign new_n9788_ = new_n7300_ & new_n7273_;
  assign new_n6973_ = ~new_n9788_;
  assign new_n9802_ = new_n9803_ & new_n7312_;
  assign new_n6974_ = ~new_n9802_;
  assign new_n9887_ = new_n7278_ & new_n7295_;
  assign new_n6975_ = ~new_n9887_;
  assign new_n9984_ = new_n7290_ & new_n7412_;
  assign new_n6976_ = ~new_n9984_;
  assign new_n6977_ = ~new_n9677_;
  assign new_n7542_ = ~new_n8820_;
  assign new_n6978_ = ~new_n8468_;
  assign new_n6979_ = ~new_n11114_;
  assign new_n6980_ = ~new_n10586_;
  assign new_n6981_ = ~new_n10005_;
  assign new_n6982_ = ~new_n10033_;
  assign new_n6983_ = ~new_n10054_;
  assign new_n6984_ = ~new_n10063_;
  assign new_n6985_ = ~new_n10042_;
  assign new_n6986_ = ~new_n10095_;
  assign new_n6987_ = ~new_n10185_;
  assign new_n7543_ = ~new_n8473_;
  assign new_n6988_ = ~new_n10195_;
  assign new_n6989_ = ~new_n10208_;
  assign new_n6990_ = ~new_n10219_;
  assign new_n6991_ = ~new_n10228_;
  assign new_n6992_ = ~new_n10241_;
  assign new_n6993_ = ~new_n10164_;
  assign new_n6994_ = ~new_n10150_;
  assign new_n11103_ = new_n9265_ & new_n11105_;
  assign new_n6995_ = ~new_n11103_;
  assign new_n10324_ = new_n7545_ & new_n7255_;
  assign new_n7544_ = ~new_n8115_;
  assign new_n6996_ = ~new_n10324_;
  assign new_n6997_ = ~new_n11381_;
  assign new_n6998_ = ~new_n11417_;
  assign new_n11294_ = new_n11434_ & new_n9537_;
  assign new_n6999_ = ~new_n11294_;
  assign new_n11447_ = new_n7481_ & new_n9338_;
  assign new_n7000_ = ~new_n11447_;
  assign new_n11432_ = new_n7468_ & new_n9494_;
  assign new_n7001_ = ~new_n11432_;
  assign new_n11428_ = new_n9532_ & new_n9530_;
  assign new_n7545_ = ~new_n7701_;
  assign new_n7002_ = ~new_n11428_;
  assign new_n7003_ = ~new_n7722_;
  assign new_n7004_ = ~new_n7819_;
  assign new_n7005_ = ~new_n7836_;
  assign new_n7006_ = ~new_n7853_;
  assign new_n7007_ = ~new_n7870_;
  assign new_n7008_ = ~new_n8551_;
  assign new_n7009_ = ~new_n7887_;
  assign new_n7010_ = ~new_n8572_;
  assign new_n7011_ = ~new_n7904_;
  assign new_n7546_ = ~new_n8629_;
  assign new_n7012_ = ~new_n7921_;
  assign new_n7013_ = ~new_n7938_;
  assign new_n7014_ = ~new_n7955_;
  assign new_n7015_ = ~new_n7972_;
  assign new_n7016_ = ~new_n7989_;
  assign new_n7017_ = ~new_n8006_;
  assign new_n7018_ = ~new_n8023_;
  assign new_n7019_ = ~new_n8040_;
  assign new_n7020_ = ~new_n8822_;
  assign new_n7021_ = ~new_n8057_;
  assign new_n7547_ = ~new_n9278_;
  assign new_n8865_ = new_n8889_ & new_n8899_;
  assign new_n7548_ = ~new_n7580_;
  assign new_n7549_ = ~new_n8274_;
  assign new_n7550_ = ~new_n9282_;
  assign new_n7074_ = ~new_n9647_;
  assign new_n7551_ = ~new_n10635_;
  assign new_n7552_ = ~new_n9313_;
  assign new_n9313_ = new_n7553_ & STATE_REG;
  assign new_n7553_ = ~new_n9311_;
  assign new_n9311_ = STATE_REG & new_n9536_;
  assign new_n7554_ = ~new_n7589_;
  assign new_n7555_ = ~new_n9551_;
  assign new_n7556_ = ~new_n9568_;
  assign new_n7557_ = ~new_n9680_;
  assign new_n7558_ = ~new_n7793_;
  assign new_n7075_ = ~new_n9725_;
  assign new_n7559_ = ~new_n7809_;
  assign new_n7809_ = new_n9269_ & new_n7772_;
  assign new_n7560_ = ~new_n8291_;
  assign new_n7561_ = ~new_n7798_;
  assign new_n7562_ = ~new_n10712_;
  assign new_n7563_ = ~new_n10713_;
  assign new_n7564_ = ~new_n8304_;
  assign new_n7565_ = ~new_n8407_;
  assign n1341 = new_n11153_ & new_n9540_;
  assign new_n7566_ = ~n1341;
  assign new_n9299_ = new_n10319_ & new_n7269_;
  assign new_n7567_ = ~new_n9293_;
  assign new_n7568_ = ~new_n7772_;
  assign new_n7569_ = ~new_n9685_;
  assign n998 = new_n6845_ | new_n6720_;
  assign new_n7579_ = new_n7548_ | new_n7189_;
  assign new_n7585_ = new_n7488_ | new_n7582_;
  assign new_n7582_ = ~new_n7354_ ^ REG2_REG_13_;
  assign new_n7584_ = new_n6311_ & new_n7554_;
  assign n994 = new_n6846_ | new_n6721_;
  assign new_n7600_ = new_n7601_ | new_n7488_;
  assign new_n7076_ = ~new_n9299_;
  assign new_n7599_ = new_n6312_ & new_n7554_;
  assign new_n7607_ = new_n7548_ | new_n7190_;
  assign new_n7601_ = ~new_n7357_ ^ REG2_REG_14_;
  assign n990 = new_n6847_ | new_n6722_;
  assign new_n7620_ = new_n7548_ | new_n7191_;
  assign new_n7625_ = new_n7622_ | new_n7488_;
  assign new_n7622_ = ~new_n7353_ ^ REG2_REG_15_;
  assign new_n7624_ = new_n6313_ & new_n7554_;
  assign n986 = new_n6848_ | new_n6723_;
  assign new_n7639_ = ~new_n7640_ ^ new_n7722_;
  assign new_n7077_ = ~new_n11268_;
  assign new_n7637_ = new_n6314_ & new_n7554_;
  assign new_n7642_ = ~new_n7493_ ^ new_n7644_;
  assign new_n7649_ = ~REG2_REG_16_ ^ new_n7493_;
  assign new_n7650_ = ~new_n7722_ ^ REG1_REG_16_;
  assign n982 = new_n6849_ | new_n6724_;
  assign new_n7661_ = ~REG2_REG_17_ ^ new_n7490_;
  assign new_n7663_ = ~REG1_REG_17_ ^ new_n7489_;
  assign new_n7668_ = ~new_n7489_ ^ new_n7669_;
  assign new_n7666_ = new_n6315_ & new_n7554_;
  assign new_n7671_ = ~new_n7490_ ^ new_n7672_;
  assign new_n11230_ = new_n11370_ & new_n7145_;
  assign n978 = new_n6850_ | new_n6725_;
  assign new_n7682_ = ~new_n7491_ ^ new_n7684_;
  assign new_n7680_ = new_n6316_ & new_n7554_;
  assign new_n7686_ = ~new_n7492_ ^ new_n7688_;
  assign new_n7693_ = ~REG2_REG_18_ ^ new_n7492_;
  assign new_n7694_ = ~REG1_REG_18_ ^ new_n7491_;
  assign n974 = new_n6851_ | new_n6726_;
  assign new_n7705_ = ~REG2_REG_19_ ^ new_n7332_;
  assign new_n7707_ = ~REG1_REG_19_ ^ new_n7331_;
  assign new_n7712_ = new_n7331_ ^ REG1_REG_19_;
  assign new_n7078_ = ~new_n11230_;
  assign new_n7684_ = ~REG1_REG_18_;
  assign new_n7715_ = new_n7537_ | new_n7491_;
  assign new_n7669_ = ~REG1_REG_17_;
  assign new_n7718_ = new_n7540_ | new_n7489_;
  assign new_n7640_ = ~REG1_REG_16_;
  assign new_n7732_ = REG1_REG_12_ & new_n7207_;
  assign new_n7729_ = new_n7734_ & new_n7304_;
  assign new_n7735_ = new_n7207_ & new_n6457_;
  assign new_n7737_ = ~REG1_REG_12_;
  assign new_n7734_ = ~REG1_REG_14_;
  assign new_n7079_ = ~new_n11171_;
  assign new_n7710_ = new_n6317_ & new_n7554_;
  assign new_n7741_ = new_n7332_ ^ REG2_REG_19_;
  assign new_n7688_ = ~REG2_REG_18_;
  assign new_n7744_ = new_n7537_ | new_n7492_;
  assign new_n7672_ = ~REG2_REG_17_;
  assign new_n7747_ = new_n7540_ | new_n7490_;
  assign new_n7644_ = ~REG2_REG_16_;
  assign new_n7750_ = new_n7513_ | new_n7493_;
  assign new_n7754_ = ~REG2_REG_15_;
  assign new_n7753_ = new_n7463_ | new_n7353_;
  assign new_n7029_ = ~new_n8179_;
  assign new_n11078_ = new_n11406_ & new_n7148_;
  assign new_n7758_ = ~REG2_REG_14_;
  assign new_n7757_ = new_n7455_ | new_n7357_;
  assign new_n7762_ = ~REG2_REG_13_;
  assign new_n7761_ = new_n7464_ | new_n7354_;
  assign new_n7765_ = new_n7505_ | new_n7510_;
  assign n969 = new_n6852_ | new_n6727_;
  assign n964 = new_n6853_ | new_n6728_;
  assign new_n7781_ = new_n7176_ & new_n7351_;
  assign n959 = new_n6854_ | new_n6729_;
  assign new_n7786_ = new_n7788_ & new_n6458_;
  assign new_n7080_ = ~new_n11078_;
  assign new_n7788_ = new_n7568_ | new_n7200_;
  assign n954 = ~new_n6013_ | ~new_n5724_;
  assign n949 = ~new_n6014_ | ~new_n5725_;
  assign n944 = ~new_n6015_ | ~new_n5726_;
  assign n939 = ~new_n6016_ | ~new_n5727_;
  assign n934 = ~new_n6017_ | ~new_n5728_;
  assign n929 = ~new_n6018_ | ~new_n5729_;
  assign n924 = ~new_n6019_ | ~new_n5730_;
  assign n919 = ~new_n6020_ | ~new_n5731_;
  assign n914 = ~new_n6021_ | ~new_n5732_;
  assign new_n8406_ = new_n7122_ & new_n7521_;
  assign n909 = ~new_n6022_ | ~new_n5733_;
  assign n904 = ~new_n6023_ | ~new_n5734_;
  assign n899 = ~new_n6024_ | ~new_n5735_;
  assign n894 = ~new_n6025_ | ~new_n5736_;
  assign n889 = ~new_n6026_ | ~new_n5737_;
  assign n884 = ~new_n6027_ | ~new_n5738_;
  assign n879 = ~new_n6028_ | ~new_n5739_;
  assign n874 = ~new_n6029_ | ~new_n5740_;
  assign n869 = ~new_n6030_ | ~new_n5741_;
  assign n864 = ~new_n6031_ | ~new_n5742_;
  assign new_n7081_ = ~new_n8406_;
  assign new_n8114_ = new_n7544_ | new_n6730_;
  assign n859 = ~new_n6032_ | ~new_n5743_;
  assign n854 = ~new_n6033_ | ~new_n5744_;
  assign new_n8150_ = new_n7544_ | new_n6731_;
  assign n849 = ~new_n6034_ | ~new_n5745_;
  assign n844 = ~new_n6035_ | ~new_n5746_;
  assign new_n8185_ = new_n7544_ | new_n6732_;
  assign n839 = ~new_n6036_ | ~new_n5747_;
  assign n834 = ~new_n6037_ | ~new_n5748_;
  assign new_n8220_ = new_n7544_ | new_n6733_;
  assign new_n8449_ = new_n8479_ & new_n8508_;
  assign new_n8217_ = new_n8223_ & new_n7558_;
  assign n829 = ~new_n6038_ | ~new_n5749_;
  assign n824 = ~new_n6039_ | ~new_n5750_;
  assign new_n8253_ = new_n7544_ | new_n6734_;
  assign n819 = ~new_n6040_ | ~new_n5751_;
  assign n814 = new_n6855_ | new_n6735_;
  assign new_n8284_ = new_n8286_ & new_n6460_;
  assign new_n8286_ = new_n7568_ | new_n6736_;
  assign new_n8289_ = new_n7560_ | new_n8292_;
  assign new_n7814_ = new_n7772_ & new_n8295_;
  assign new_n7082_ = ~new_n8449_;
  assign n809 = ~new_n6041_ | ~new_n5752_;
  assign n804 = ~new_n6042_ | ~new_n5753_;
  assign n799 = ~new_n6043_ | ~new_n5754_;
  assign n794 = ~new_n6044_ | ~new_n5755_;
  assign n789 = ~new_n6045_ | ~new_n5756_;
  assign n784 = ~new_n6046_ | ~new_n5757_;
  assign n779 = ~new_n6047_ | ~new_n5758_;
  assign n774 = ~new_n6048_ | ~new_n5759_;
  assign n769 = ~new_n6049_ | ~new_n5760_;
  assign n764 = ~new_n6050_ | ~new_n5761_;
  assign new_n8508_ = new_n8542_ & new_n8569_;
  assign n759 = ~new_n6051_ | ~new_n5762_;
  assign n754 = ~new_n6052_ | ~new_n5763_;
  assign n749 = ~new_n6053_ | ~new_n5764_;
  assign n744 = ~new_n6054_ | ~new_n5765_;
  assign n739 = ~new_n6055_ | ~new_n5766_;
  assign n734 = ~new_n6056_ | ~new_n5767_;
  assign n729 = ~new_n6057_ | ~new_n5768_;
  assign n724 = ~new_n6058_ | ~new_n5769_;
  assign n719 = ~new_n6059_ | ~new_n5770_;
  assign n714 = ~new_n6060_ | ~new_n5771_;
  assign new_n7083_ = ~new_n8508_;
  assign n709 = ~new_n6061_ | ~new_n5772_;
  assign n704 = ~new_n6062_ | ~new_n5773_;
  assign n699 = ~new_n6063_ | ~new_n5774_;
  assign n694 = ~new_n6064_ | ~new_n5775_;
  assign n689 = ~new_n6065_ | ~new_n5776_;
  assign n684 = ~new_n6066_ | ~new_n5777_;
  assign n679 = ~new_n6067_ | ~new_n5778_;
  assign n674 = ~new_n6068_ | ~new_n5779_;
  assign n669 = ~new_n6069_ | ~new_n5780_;
  assign n664 = ~new_n6070_ | ~new_n5781_;
  assign new_n8569_ = new_n8592_ & new_n8634_;
  assign n659 = ~new_n6071_ | ~new_n5782_;
  assign n654 = ~new_n6072_ | ~new_n5783_;
  assign n649 = ~new_n6073_ | ~new_n5784_;
  assign new_n8402_ = new_n6318_ & new_n7081_;
  assign new_n7775_ = ~new_n7351_ ^ new_n7431_;
  assign n644 = ~new_n6074_ | ~new_n5785_;
  assign new_n8414_ = new_n7461_ & new_n7407_;
  assign n639 = ~new_n6076_ | ~new_n5786_;
  assign new_n8310_ = new_n6856_ | new_n6737_;
  assign new_n7799_ = ~new_n8449_ ^ new_n8415_;
  assign new_n7084_ = ~new_n8569_;
  assign new_n7794_ = ~new_n6944_ ^ new_n7352_;
  assign new_n8455_ = new_n7519_ | new_n7367_;
  assign n634 = ~new_n6077_ | ~new_n5787_;
  assign new_n8313_ = new_n6857_ | new_n6738_;
  assign new_n8466_ = new_n7344_ ^ new_n8467_;
  assign new_n8470_ = new_n7462_ & new_n7543_;
  assign new_n7806_ = new_n6319_ & new_n7082_;
  assign new_n8479_ = new_n7519_ & new_n7457_;
  assign new_n7807_ = new_n7367_ ^ new_n8467_;
  assign new_n8481_ = new_n7361_ | new_n7828_;
  assign new_n7030_ = ~new_n8197_;
  assign new_n8634_ = new_n8658_ & new_n8690_;
  assign n629 = ~new_n6079_ | ~new_n5789_;
  assign new_n8316_ = new_n6859_ | new_n6739_;
  assign new_n8491_ = new_n6321_ & new_n8494_;
  assign new_n8494_ = new_n6858_ | new_n6740_;
  assign new_n8498_ = new_n7435_ & new_n7543_;
  assign new_n8501_ = new_n6320_ & new_n7091_;
  assign new_n7826_ = ~new_n8508_ ^ new_n7828_;
  assign new_n7827_ = ~new_n7361_ ^ new_n8503_;
  assign new_n8511_ = new_n7178_ & new_n8572_;
  assign new_n8516_ = new_n7177_ & new_n6465_;
  assign new_n7085_ = ~new_n8634_;
  assign n624 = ~new_n6080_ | ~new_n5790_;
  assign new_n8319_ = new_n6860_ | new_n6741_;
  assign new_n8531_ = new_n7435_ ^ new_n8532_;
  assign new_n7843_ = new_n6322_ & new_n7083_;
  assign new_n8542_ = new_n7512_ & new_n7447_;
  assign new_n7844_ = new_n8544_ & new_n6468_;
  assign new_n8546_ = new_n7298_ & new_n6469_;
  assign new_n8544_ = new_n7292_ | new_n6742_;
  assign n619 = ~new_n6082_ | ~new_n5791_;
  assign new_n8322_ = new_n6861_ | new_n6743_;
  assign new_n7086_ = ~new_n8690_;
  assign new_n8563_ = ~new_n8564_ ^ new_n8536_;
  assign new_n7860_ = ~new_n8569_ ^ new_n7862_;
  assign new_n7861_ = ~new_n8551_ ^ new_n8564_;
  assign n614 = ~new_n6083_ | ~new_n5792_;
  assign new_n8325_ = new_n6862_ | new_n6744_;
  assign new_n8582_ = new_n8583_ ^ new_n8584_;
  assign new_n8583_ = new_n7205_ | new_n8586_;
  assign new_n7877_ = new_n6323_ & new_n7084_;
  assign new_n8592_ = new_n7454_ & new_n7538_;
  assign new_n7878_ = ~new_n8572_ ^ new_n8584_;
  assign new_n7087_ = ~new_n8747_;
  assign new_n8597_ = new_n7538_ | new_n7358_;
  assign n609 = ~new_n6085_ | ~new_n5793_;
  assign new_n8328_ = new_n6864_ | new_n6745_;
  assign new_n8608_ = new_n6863_ | new_n6746_;
  assign new_n8611_ = new_n7530_ | new_n7434_;
  assign new_n8625_ = new_n7482_ & new_n7546_;
  assign new_n7894_ = ~new_n8634_ ^ new_n7896_;
  assign new_n7895_ = ~new_n7358_ ^ new_n7434_;
  assign new_n8635_ = new_n7362_ | new_n7913_;
  assign n604 = ~new_n6086_ | ~new_n5795_;
  assign new_n7088_ = ~new_n8794_;
  assign new_n8331_ = new_n6865_ | new_n6747_;
  assign new_n8649_ = new_n7226_ ^ new_n8650_;
  assign new_n7911_ = new_n6324_ & new_n7085_;
  assign new_n8658_ = new_n7509_ & new_n7395_;
  assign new_n7912_ = ~new_n7362_ ^ new_n8650_;
  assign new_n8664_ = new_n7179_ & new_n7335_;
  assign new_n8668_ = new_n6866_ | new_n7330_;
  assign new_n8665_ = new_n8673_ & new_n7166_;
  assign n599 = ~new_n6088_ | ~new_n5796_;
  assign new_n8334_ = new_n6867_ | new_n6748_;
  assign new_n7089_ = ~new_n8862_;
  assign new_n8684_ = ~new_n8652_ ^ new_n7347_;
  assign new_n8652_ = new_n7310_ | new_n8627_;
  assign new_n7928_ = ~new_n8690_ ^ new_n7930_;
  assign new_n8693_ = new_n8694_ | new_n7330_;
  assign new_n8694_ = new_n8731_ & new_n8673_;
  assign n594 = ~new_n6089_ | ~new_n5797_;
  assign new_n8337_ = new_n6868_ | new_n6749_;
  assign new_n8708_ = new_n6955_ ^ new_n8710_;
  assign new_n7945_ = new_n6325_ & new_n7086_;
  assign new_n8724_ = new_n6326_ & new_n7270_;
  assign new_n7090_ = ~new_n8916_;
  assign new_n8673_ = new_n7160_ & new_n7167_;
  assign new_n8727_ = new_n6327_ & new_n7152_;
  assign n589 = ~new_n6090_ | ~new_n5798_;
  assign new_n8340_ = new_n6869_ | new_n6750_;
  assign new_n8741_ = new_n7365_ ^ new_n8742_;
  assign new_n7962_ = ~new_n8747_ ^ new_n7964_;
  assign new_n7963_ = ~new_n8731_ ^ new_n8742_;
  assign n584 = ~new_n6092_ | ~new_n5800_;
  assign new_n8343_ = new_n6870_ | new_n6751_;
  assign new_n8760_ = new_n7225_ ^ new_n8762_;
  assign new_n8503_ = new_n7462_ & new_n7413_;
  assign new_n7979_ = new_n6328_ & new_n7087_;
  assign new_n7980_ = ~new_n7335_ ^ new_n8762_;
  assign new_n8775_ = new_n7419_ | new_n7536_;
  assign new_n8770_ = new_n7217_ | new_n8800_;
  assign n579 = ~new_n6093_ | ~new_n5802_;
  assign new_n8346_ = new_n6871_ | new_n6752_;
  assign new_n8787_ = ~new_n7223_ ^ new_n7224_;
  assign new_n7996_ = ~new_n8794_ ^ new_n7998_;
  assign new_n7997_ = new_n8795_ & new_n6491_;
  assign new_n8797_ = new_n6329_ & new_n7419_;
  assign new_n7091_ = ~new_n8503_;
  assign new_n8795_ = new_n7217_ | new_n6753_;
  assign n574 = ~new_n6098_ | ~new_n5803_;
  assign new_n8349_ = new_n6872_ | new_n6754_;
  assign new_n8013_ = new_n6330_ & new_n7088_;
  assign new_n8014_ = ~new_n7333_ ^ new_n8824_;
  assign new_n8834_ = new_n7311_ | new_n7532_;
  assign new_n8838_ = new_n6331_ & new_n7282_;
  assign n569 = ~new_n6099_ | ~new_n5804_;
  assign new_n8352_ = new_n6873_ | new_n6755_;
  assign new_n8852_ = ~new_n8822_ ^ new_n8853_;
  assign new_n10810_ = new_n10820_ & REG3_REG_20_;
  assign new_n8030_ = ~new_n8862_ ^ new_n8032_;
  assign new_n8031_ = ~new_n6945_ ^ new_n8853_;
  assign n564 = ~new_n6100_ | ~new_n5806_;
  assign new_n8355_ = new_n6874_ | new_n6756_;
  assign new_n8879_ = new_n7356_ ^ new_n8880_;
  assign new_n8047_ = new_n6332_ & new_n7089_;
  assign new_n8048_ = ~new_n6946_ ^ new_n8880_;
  assign new_n8889_ = new_n7116_ & new_n7336_;
  assign new_n8894_ = new_n7180_ & new_n6500_;
  assign new_n8898_ = new_n8952_ & new_n8899_;
endmodule



module wf_8x6 #(parameter N = 16, parameter stages = 6) ( // TOKEN_WF_MODNAME
    input [N-1:0] IN,
    input [N*stages/2-1:0] K0,
    input [N*stages/2-1:0] K1,
    input [N*stages/2-1:0] K2,
    output [N-1:0] OUT
);
    wire [N-1:0] cln_out;
    wire [N-1:0] inverted_in;
    wire [N-1:0] unpermuted_out;

//    assign inverted_in[0]  =   IN[0];
//    assign inverted_in[1]  =  !IN[1];
//    assign inverted_in[2]  =   IN[2];
//    assign inverted_in[3]  =  !IN[3];
    // TOKEN_BEGIN_INVERSIONS
    assign inverted_in[0] =  IN[0];
    assign inverted_in[1] =  IN[1];
    assign inverted_in[2] =  IN[2];
    assign inverted_in[3] = !IN[3];
    assign inverted_in[4] =  IN[4];
    assign inverted_in[5] = !IN[5];
    assign inverted_in[6] = !IN[6];
    assign inverted_in[7] =  IN[7];
    assign inverted_in[8] =  IN[8];
    assign inverted_in[9] = !IN[9];
    assign inverted_in[10] =  IN[10];
    assign inverted_in[11] =  IN[11];
    assign inverted_in[12] = !IN[12];
    assign inverted_in[13] = !IN[13];
    assign inverted_in[14] =  IN[14];
    assign inverted_in[15] = !IN[15];


    cln #(.N(N), .stages(stages)) wf_cln(
        .IN(inverted_in),
        .K0(K0),
        .K1(K1),
        .K2(K2),
        .OUT(cln_out)
    );

    assign unpermuted_out = {
//        cln_out[2],
//        cln_out[1],
//        cln_out[0],
//        cln_out[3]
        // TOKEN_BEGIN_PERMUTATION
        cln_out[14],
        cln_out[0],
        cln_out[8],
        cln_out[13],
        cln_out[3],
        cln_out[12],
        cln_out[11],
        cln_out[10],
        cln_out[15],
        cln_out[9],
        cln_out[6],
        cln_out[4],
        cln_out[2],
        cln_out[1],
        cln_out[7],
        cln_out[5]
    };


//    lut1 lut_0 (
//        .inputs(unpermuted_out[0]),
//        .outputs(OUT[0])
//    );
//
//    lut3 lut_1 (
//        .inputs(unpermuted_out[3:1]),
//        .outputs(OUT[3:1])
//    );
    // TOKEN_BEGIN_LUTS
    lut2 lut_0 (
        .inputs(unpermuted_out[1:0]),
        .outputs(OUT[1:0])
    );

    lut2 lut_1 (
        .inputs(unpermuted_out[3:2]),
        .outputs(OUT[3:2])
    );

    lut2 lut_2 (
        .inputs(unpermuted_out[5:4]),
        .outputs(OUT[5:4])
    );

    lut2 lut_3 (
        .inputs(unpermuted_out[7:6]),
        .outputs(OUT[7:6])
    );

    lut2 lut_4 (
        .inputs(unpermuted_out[9:8]),
        .outputs(OUT[9:8])
    );

    lut2 lut_5 (
        .inputs(unpermuted_out[11:10]),
        .outputs(OUT[11:10])
    );

    lut2 lut_6 (
        .inputs(unpermuted_out[13:12]),
        .outputs(OUT[13:12])
    );

    lut2 lut_7 (
        .inputs(unpermuted_out[15:14]),
        .outputs(OUT[15:14])
    );



endmodule
